//: version "1.8.7"

module jump(SignXtended, dir, PCNext, jump, PCSrc, inm26);
//: interface  /sz:(121, 80) /bd:[ Ti0>jump(74/121) Li0>PCNext[31:0](51/80) Li1>inm26[25:0](19/80) Bi0>PCSrc(85/121) Bi1>SignXtended[31:0](37/121) Ro0<dir[31:0](36/80) ]
input jump;    //: /sn:0 {0}(503,158)(503,124){1}
input PCSrc;    //: /sn:0 /dp:1 {0}(433,134)(433,180){1}
input [25:0] inm26;    //: /sn:0 {0}(139,76)(272,76){1}
supply0 w3;    //: /sn:0 {0}(328,47)(328,97){1}
output [31:0] dir;    //: /sn:0 /dp:1 {0}(516,101)(568,101){1}
input [31:0] PCNext;    //: /sn:0 /dp:1 {0}(417,101)(353,101)(353,83)(301,83)(301,103){1}
//: {2}(303,105)(314,105){3}
//: {4}(299,105)(203,105){5}
//: {6}(202,105)(139,105){7}
input [31:0] SignXtended;    //: /sn:0 /dp:1 {0}(314,137)(292,137)(292,175){1}
wire w6;    //: /sn:0 /dp:1 {0}(328,145)(328,155){1}
wire [31:0] w7;    //: /sn:0 {0}(417,121)(343,121){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(487,111)(446,111){1}
wire [5:0] w1;    //: /sn:0 {0}(203,100)(203,66)(272,66){1}
wire [31:0] w2;    //: /sn:0 {0}(278,71)(461,71)(461,91)(487,91){1}
//: enddecls

  concat g4 (.I0(inm26), .I1(w1), .Z(w2));   //: @(277,71) /sn:0 /w:[ 1 1 0 ] /dr:0
  mux g8 (.I0(PCNext), .I1(w7), .S(PCSrc), .Z(w0));   //: @(433,111) /sn:0 /R:1 /w:[ 0 0 0 1 ] /ss:0 /do:1
  //: input g3 (SignXtended) @(292,177) /sn:0 /R:1 /w:[ 1 ]
  //: output g2 (dir) @(565,101) /sn:0 /w:[ 1 ]
  //: input g1 (PCNext) @(137,105) /sn:0 /w:[ 7 ]
  //: joint g10 (PCNext) @(301, 105) /w:[ 2 1 4 -1 ]
  add g6 (.A(SignXtended), .B(PCNext), .S(w7), .CI(w3), .CO(w6));   //: @(330,121) /sn:0 /R:1 /w:[ 0 3 1 1 0 ]
  mux g7 (.I0(w0), .I1(w2), .S(jump), .Z(dir));   //: @(503,101) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:0 /do:0
  //: input g9 (jump) @(503,160) /sn:0 /R:1 /w:[ 0 ]
  //: supply0 g12 (w3) @(328,41) /sn:0 /R:2 /w:[ 0 ]
  tran g5(.Z(w1), .I(PCNext[31:26]));   //: @(203,103) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:0
  //: input g11 (PCSrc) @(433,182) /sn:0 /R:1 /w:[ 1 ]
  //: input g0 (inm26) @(137,76) /sn:0 /w:[ 0 ]

endmodule

module memoria(RD, WD, Addr, MemRead, MemWrite, clk);
//: interface  /sz:(297, 200) /bd:[ Ti0>MemWrite(147/297) Li0>WD[31:0](133/200) Li1>Addr[31:0](37/200) Bi0>clk(224/297) Bi1>MemRead(133/297) Ro0<RD[31:0](82/200) ]
supply0 w0;    //: /sn:0 {0}(715,297)(715,278){1}
input [31:0] Addr;    //: /sn:0 {0}(668,253)(704,253){1}
input [31:0] WD;    //: /sn:0 /dp:1 {0}(786,224)(786,201)(771,201){1}
input MemWrite;    //: /sn:0 {0}(623,163)(718,163){1}
//: {2}(722,163)(809,163)(809,232)(791,232){3}
//: {4}(720,165)(720,181){5}
input clk;    //: /sn:0 {0}(637,147)(725,147)(725,181){1}
output [31:0] RD;    //: /sn:0 {0}(833,251)(788,251){1}
//: {2}(786,249)(786,240){3}
//: {4}(784,251)(739,251){5}
input MemRead;    //: /sn:0 {0}(683,339)(729,339)(729,278){1}
wire w9;    //: /sn:0 {0}(722,202)(722,228){1}
//: enddecls

  //: output g4 (RD) @(830,251) /sn:0 /w:[ 0 ]
  bufif1 g8 (.Z(RD), .I(WD), .E(MemWrite));   //: @(786,230) /sn:0 /R:3 /w:[ 3 0 3 ]
  //: input g3 (WD) @(769,201) /sn:0 /w:[ 1 ]
  //: supply0 g2 (w0) @(715,303) /sn:0 /w:[ 0 ]
  //: input g1 (Addr) @(666,253) /sn:0 /w:[ 0 ]
  //: joint g10 (MemWrite) @(720, 163) /w:[ 2 -1 1 4 ]
  //: input g6 (MemRead) @(681,339) /sn:0 /w:[ 0 ]
  //: input g7 (MemWrite) @(621,163) /sn:0 /w:[ 0 ]
  nand g9 (.I0(clk), .I1(MemWrite), .Z(w9));   //: @(722,192) /sn:0 /R:3 /w:[ 1 5 0 ]
  //: input g5 (clk) @(635,147) /sn:0 /w:[ 0 ]
  //: joint g11 (RD) @(786, 251) /w:[ 1 2 4 -1 ]
  ram g0 (.A(Addr), .D(RD), .WE(w9), .OE(!MemRead), .CS(w0));   //: @(722,252) /sn:0 /w:[ 1 5 1 1 1 ]

endmodule

module ALU(AluOp, Z, B, AluResult, A);
//: interface  /sz:(40, 40) /bd:[ Ti0>op[3:0](20/40) Li0>a[31:0](10/40) Li1>b[31:0](30/40) Ro0<Q[31:0](30/40) Ro1<Z(10/40) ]
input [31:0] B;    //: /sn:0 /dp:1 {0}(626,444)(575,444)(575,381){1}
//: {2}(577,379)(695,379)(695,443)(740,443){3}
//: {4}(575,377)(575,285)(483,285){5}
input [31:0] A;    //: /sn:0 /dp:8 {0}(792,239)(727,239){1}
//: {2}(723,239)(663,239){3}
//: {4}(659,239)(529,239)(529,226)(483,226){5}
//: {6}(661,241)(661,318)(919,318){7}
//: {8}(725,241)(725,288)(801,288){9}
output Z;    //: /sn:0 /dp:1 {0}(1393,261)(1328,261){1}
supply0 [30:0] w12;    //: /sn:0 {0}(1000,349)(1000,372)(1001,372){1}
output [31:0] AluResult;    //: /sn:0 {0}(1307,261)(1234,261)(1234,290){1}
//: {2}(1232,292)(1180,292)(1180,294)(1130,294){3}
//: {4}(1234,294)(1234,327)(1350,327){5}
input [3:0] AluOp;    //: /sn:0 {0}(510,533)(755,533){1}
//: {2}(756,533)(1114,533){3}
//: {4}(1115,533)(1169,533){5}
wire [1:0] w4;    //: /sn:0 {0}(1115,528)(1115,521)(1117,521)(1117,317){1}
wire w0;    //: /sn:0 {0}(968,338)(968,382)(1001,382){1}
wire [31:0] w3;    //: /sn:0 {0}(642,444)(671,444)(671,423)(740,423){1}
wire [31:0] w10;    //: /sn:0 {0}(948,334)(967,334){1}
//: {2}(968,334)(990,334)(990,300)(1101,300){3}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(1101,288)(875,288)(875,286)(822,286){1}
wire [31:0] w8;    //: /sn:0 /dp:1 {0}(919,350)(905,350)(905,433)(793,433){1}
//: {2}(791,431)(791,399){3}
//: {4}(791,395)(791,244)(792,244){5}
//: {6}(789,397)(761,397)(761,283)(801,283){7}
//: {8}(789,433)(769,433){9}
wire [31:0] w2;    //: /sn:0 {0}(813,242)(1091,242)(1091,276)(1101,276){1}
wire w11;    //: /sn:0 /dp:1 {0}(933,391)(933,358){1}
wire w5;    //: /sn:0 {0}(756,528)(756,491){1}
//: {2}(758,489)(847,489)(847,300)(933,300)(933,310){3}
//: {4}(756,487)(756,456){5}
wire [31:0] w9;    //: /sn:0 /dp:1 {0}(1007,377)(1110,377)(1110,327)(1091,327)(1091,312)(1101,312){1}
//: enddecls

  not g4 (.I(B), .Z(w3));   //: @(632,444) /sn:0 /w:[ 0 0 ]
  tran g8(.Z(w5), .I(AluOp[2]));   //: @(756,531) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  mux g16 (.I0(w2), .I1(w1), .I2(w10), .I3(w9), .S(w4), .Z(AluResult));   //: @(1117,294) /sn:0 /R:1 /w:[ 1 0 3 1 1 3 ] /ss:0 /do:1
  and g3 (.I0(A), .I1(w8), .Z(w2));   //: @(803,242) /sn:0 /w:[ 0 5 0 ]
  concat g17 (.I0(w0), .I1(w12), .Z(w9));   //: @(1006,377) /sn:0 /w:[ 1 1 0 ] /dr:0
  //: input g2 (AluOp) @(508,533) /sn:0 /w:[ 0 ]
  //: joint g23 (AluResult) @(1234, 292) /w:[ -1 1 2 4 ]
  //: output g24 (Z) @(1390,261) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(481,285) /sn:0 /w:[ 5 ]
  tran g18(.Z(w0), .I(w10[31]));   //: @(968,332) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g10 (w5) @(756, 489) /w:[ 2 4 -1 1 ]
  //: joint g6 (B) @(575, 379) /w:[ 2 4 -1 1 ]
  or g7 (.I0(w8), .I1(A), .Z(w1));   //: @(812,286) /sn:0 /w:[ 7 9 1 ]
  add g9 (.A(w8), .B(A), .S(w10), .CI(w5), .CO(w11));   //: @(935,334) /sn:0 /R:1 /w:[ 0 7 0 3 1 ]
  //: output g22 (AluResult) @(1347,327) /sn:0 /w:[ 5 ]
  //: joint g12 (A) @(661, 239) /w:[ 3 -1 4 6 ]
  //: joint g14 (w8) @(791, 433) /w:[ 1 2 8 -1 ]
  mux g5 (.I0(B), .I1(w3), .S(w5), .Z(w8));   //: @(756,433) /sn:0 /R:1 /w:[ 3 1 5 9 ] /ss:0 /do:0
  led g11 (.I(w11));   //: @(933,398) /sn:0 /R:2 /w:[ 0 ] /type:0
  nor g21 (.I0(AluResult), .Z(Z));   //: @(1318,261) /sn:0 /w:[ 0 1 ]
  //: supply0 g19 (w12) @(1000,343) /sn:0 /R:2 /w:[ 0 ]
  tran g20(.Z(w4), .I(AluOp[1:0]));   //: @(1115,531) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:0
  //: joint g15 (w8) @(791, 397) /w:[ -1 4 6 3 ]
  //: input g0 (A) @(481,226) /sn:0 /w:[ 5 ]
  //: joint g13 (A) @(725, 239) /w:[ 1 -1 2 8 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Li0>Read1[4:0](32/182) Li1>Read2[4:0](72/182) Li2>Write[4:0](108/182) Li3>WriteData[31:0](148/182) Bi0>clk(108/147) Bi1>RegWrite(40/147) Ro0<Data1[31:0](47/182) Ro1<Data2[31:0](139/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clk, clr, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Li0>clk(59/69) Li1>RegWr(47/69) Li2>SB[2:0](22/69) Li3>SA[2:0](11/69) Li4>SD[2:0](35/69) Ri0>clr(35/69) Bo0<BOUT[31:0](65/98) Bo1<AOUT[31:0](37/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module Fetch(Inst, Reset, Clk, PCIn, PCOut);
//: interface  /sz:(107, 96) /bd:[ Ti0>PCIn[31:0](76/107) Ti1>PCIn[31:0](76/107) Li0>Clk(65/96) Li1>Reset(22/96) Li2>Reset(22/96) Li3>Clk(65/96) To0<PCOut[31:0](28/107) To1<PCOut[31:0](28/107) Ro0<Inst[31:0](49/96) Ro1<Inst[31:0](49/96) ]
supply0 w13;    //: /sn:0 {0}(348,222)(348,195){1}
output [31:0] PCOut;    //: /sn:0 /dp:1 {0}(429,76)(482,76){1}
input Clk;    //: /sn:0 {0}(188,208)(238,208)(238,185){1}
output [31:0] Inst;    //: /sn:0 {0}(427,168)(365,168){1}
input [31:0] PCIn;    //: /sn:0 {0}(148,147)(227,147){1}
input Reset;    //: /sn:0 {0}(182,91)(233,91)(233,109){1}
supply0 w14;    //: /sn:0 {0}(258,73)(258,99)(243,99)(243,109){1}
supply0 w15;    //: /sn:0 {0}(439,39)(414,39)(414,52){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(352,46)(352,60)(400,60){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(248,147)(301,147){1}
//: {2}(305,147)(326,147)(326,170)(330,170){3}
//: {4}(303,145)(303,92)(400,92){5}
wire w12;    //: /sn:0 {0}(414,100)(414,110){1}
//: enddecls

  //: output g8 (Inst) @(424,168) /sn:0 /w:[ 0 ]
  //: supply0 g4 (w14) @(258,67) /sn:0 /R:2 /w:[ 0 ]
  //: supply0 g3 (w13) @(348,228) /sn:0 /w:[ 0 ]
  add g2 (.A(w3), .B(w0), .S(PCOut), .CI(w15), .CO(w12));   //: @(416,76) /sn:0 /R:1 /w:[ 5 1 0 1 0 ]
  register g1 (.Q(w3), .D(PCIn), .EN(w14), .CLR(!Reset), .CK(Clk));   //: @(238,147) /sn:0 /R:1 /w:[ 0 1 1 1 1 ]
  //: input g10 (Reset) @(180,91) /sn:0 /w:[ 0 ]
  //: joint g6 (w3) @(303, 147) /w:[ 2 4 1 -1 ]
  //: input g9 (Clk) @(186,208) /sn:0 /w:[ 0 ]
  //: dip g7 (w0) @(352,36) /sn:0 /w:[ 0 ] /st:1
  //: input g12 (PCIn) @(146,147) /sn:0 /w:[ 0 ]
  //: supply0 g5 (w15) @(445,39) /sn:0 /R:1 /w:[ 0 ]
  //: output g11 (PCOut) @(479,76) /sn:0 /w:[ 1 ]
  rom g0 (.A(w3), .D(Inst), .OE(w13));   //: @(348,169) /sn:0 /w:[ 3 1 1 ] /mem:"/media/sf_Carpeta_Compartida_Linux/EC-2/mult.mem"

endmodule

module main;    //: root_module
wire [31:0] w13;    //: /sn:0 {0}(956,271)(977,271){1}
//: {2}(981,271)(1001,271){3}
//: {4}(979,269)(979,246)(989,246)(989,198)(1143,198)(1143,180){5}
//: {6}(979,273)(979,400)(1211,400)(1211,319)(1256,319){7}
wire [4:0] w16;    //: /sn:0 {0}(548,200)(486,200){1}
wire w6;    //: /sn:0 {0}(1079,218)(1094,218)(1094,248){1}
wire w7;    //: /sn:0 {0}(796,-4)(808,-4)(808,13){1}
wire [25:0] w4;    //: /sn:0 {0}(733,33)(486,33){1}
wire [31:0] w25;    //: /sn:0 {0}(712,340)(771,340)(771,283){1}
//: {2}(773,281)(801,281){3}
//: {4}(771,279)(771,95){5}
wire [31:0] w22;    //: /sn:0 /dp:1 {0}(830,271)(884,271){1}
wire [31:0] w0;    //: /sn:0 {0}(393,352)(393,-20)(879,-20)(879,28){1}
//: {2}(881,30)(1054,30)(1054,22){3}
//: {4}(879,32)(879,50)(856,50){5}
wire [15:0] w20;    //: /sn:0 {0}(548,335)(486,335){1}
wire w18;    //: /sn:0 {0}(613,108)(634,108)(634,134){1}
wire w19;    //: /sn:0 {0}(1258,247)(1272,247)(1272,286){1}
wire [3:0] w12;    //: /sn:0 {0}(920,163)(920,222){1}
wire w10;    //: /sn:0 {0}(526,257)(548,257){1}
wire [31:0] w23;    //: /sn:0 {0}(1256,299)(1189,299){1}
wire w21;    //: /sn:0 /dp:1 {0}(974,225)(974,239)(956,239){1}
wire [31:0] w24;    //: /sn:0 {0}(1001,330)(743,330)(743,263){1}
//: {2}(745,261)(778,261){3}
//: {4}(782,261)(801,261){5}
//: {6}(780,263)(780,386){7}
//: {8}(741,261)(712,261){9}
wire w1;    //: /sn:0 {0}(654,540)(660,540)(660,380){1}
wire [31:0] w31;    //: /sn:0 /dp:1 {0}(1285,309)(1293,309)(1293,366){1}
//: {2}(1295,368)(1421,368)(1421,342){3}
//: {4}(1293,370)(1293,433)(534,433)(534,288)(548,288){5}
wire [31:0] w8;    //: /sn:0 {0}(482,25)(482,32){1}
//: {2}(482,33)(482,168){3}
//: {4}(482,169)(482,199){5}
//: {6}(482,200)(482,231){7}
//: {8}(482,232)(482,295){9}
//: {10}(480,297)(207,297)(207,257){11}
//: {12}(482,299)(482,334){13}
//: {14}(482,335)(482,402)(425,402){15}
wire [4:0] w17;    //: /sn:0 {0}(548,232)(486,232){1}
wire w28;    //: /sn:0 {0}(1142,372)(1142,569)(606,569){1}
//: {2}(604,567)(604,380){3}
//: {4}(602,569)(278,569){5}
//: {6}(276,567)(276,418)(316,418){7}
//: {8}(274,569)(166,569){9}
wire w14;    //: /sn:0 {0}(810,213)(817,213)(817,248){1}
wire w2;    //: /sn:0 {0}(268,375)(316,375){1}
wire [31:0] w11;    //: /sn:0 {0}(884,239)(843,239)(843,186){1}
//: {2}(845,184)(1001,184)(1001,127){3}
//: {4}(841,184)(712,184){5}
wire [4:0] w15;    //: /sn:0 {0}(548,169)(486,169){1}
wire w5;    //: /sn:0 {0}(1073,454)(1085,454)(1085,372){1}
wire [31:0] w26;    //: /sn:0 {0}(345,352)(345,65)(733,65){1}
wire w9;    //: /sn:0 {0}(811,133)(819,133)(819,95){1}
//: enddecls

  clock g4 (.Z(w28));   //: @(153,569) /sn:0 /w:[ 9 ] /omega:2000 /phi:0 /duty:50
  tran g8(.Z(w15), .I(w8[25:21]));   //: @(480,169) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  //: switch g16 (w18) @(596,108) /sn:0 /w:[ 0 ] /st:0
  Read g3 (.RegWrite(w18), .SignExIn(w20), .WriteData(w31), .RegDst(w10), .WR(w17), .R2(w16), .R1(w15), .clr(w1), .clk(w28), .SignExOut(w25), .RD2(w24), .RD1(w11));   //: @(549, 135) /sz:(162, 244) /sn:0 /p:[ Ti0>1 Li0>0 Li1>5 Li2>1 Li3>0 Li4>0 Li5>0 Bi0>1 Bi1>3 Ro0<0 Ro1<9 Ro2<5 ]
  //: switch g17 (w14) @(793,213) /sn:0 /w:[ 0 ] /st:0
  //: switch g26 (w19) @(1241,247) /sn:0 /w:[ 0 ] /st:0
  ALU g2 (.AluOp(w12), .A(w11), .B(w22), .AluResult(w13), .Z(w21));   //: @(885, 223) /sz:(70, 65) /sn:0 /p:[ Ti0>1 Li0>0 Li1>1 Ro0<0 Ro1<1 ]
  //: joint g23 (w13) @(979, 271) /w:[ 2 4 1 6 ]
  led g30 (.I(w0));   //: @(1054,15) /sn:0 /w:[ 3 ] /type:2
  jump g1 (.jump(w7), .PCNext(w26), .inm26(w4), .PCSrc(w9), .SignXtended(w25), .dir(w0));   //: @(734, 14) /sz:(121, 80) /sn:0 /p:[ Ti0>1 Li0>1 Li1>0 Bi0>1 Bi1>5 Ro0<5 ]
  //: switch g24 (w5) @(1056,454) /sn:0 /w:[ 0 ] /st:0
  //: joint g39 (w24) @(780, 261) /w:[ 4 -1 3 6 ]
  //: joint g29 (w31) @(1293, 368) /w:[ 2 1 -1 4 ]
  led g18 (.I(w21));   //: @(974,218) /sn:0 /w:[ 0 ] /type:0
  tran g10(.Z(w17), .I(w8[15:11]));   //: @(480,232) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: switch g25 (w6) @(1062,218) /sn:0 /w:[ 0 ] /st:0
  //: switch g6 (w2) @(251,375) /sn:0 /w:[ 0 ] /st:0
  //: switch g7 (w1) @(637,540) /sn:0 /w:[ 0 ] /st:0
  tran g9(.Z(w16), .I(w8[20:16]));   //: @(480,200) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  //: switch g35 (w7) @(779,-4) /sn:0 /w:[ 0 ] /st:0
  //: joint g22 (w28) @(604, 569) /w:[ 1 2 4 -1 ]
  //: joint g31 (w0) @(879, 30) /w:[ 2 1 -1 4 ]
  //: joint g33 (w8) @(482, 297) /w:[ -1 9 10 12 ]
  led g36 (.I(w11));   //: @(1001,120) /sn:0 /w:[ 3 ] /type:2
  led g40 (.I(w13));   //: @(1143,173) /sn:0 /w:[ 5 ] /type:2
  tran g12(.Z(w4), .I(w8[25:0]));   //: @(480,33) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  led g28 (.I(w31));   //: @(1421,335) /sn:0 /w:[ 3 ] /type:2
  //: switch g34 (w9) @(794,133) /sn:0 /w:[ 0 ] /st:0
  //: joint g14 (w25) @(771, 281) /w:[ 2 4 -1 1 ]
  //: joint g5 (w28) @(276, 569) /w:[ 5 6 8 -1 ]
  tran g11(.Z(w20), .I(w8[15:0]));   //: @(480,335) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  memoria g19 (.MemWrite(w6), .WD(w24), .Addr(w13), .clk(w28), .MemRead(w5), .RD(w23));   //: @(1002, 249) /sz:(186, 122) /sn:0 /p:[ Ti0>1 Li0>0 Li1>3 Bi0>0 Bi1>1 Ro0<1 ]
  mux g21 (.I0(w13), .I1(w23), .S(w19), .Z(w31));   //: @(1272,309) /sn:0 /R:1 /w:[ 7 0 1 0 ] /ss:1 /do:0
  //: joint g20 (w24) @(743, 261) /w:[ 2 -1 8 1 ]
  led g32 (.I(w8));   //: @(207,250) /sn:0 /w:[ 11 ] /type:2
  //: switch g15 (w10) @(509,257) /sn:0 /w:[ 0 ] /st:0
  Fetch g0 (.PCIn(w0), .Reset(w2), .Clk(w28), .PCOut(w26), .Inst(w8));   //: @(317, 353) /sz:(107, 96) /sn:0 /p:[ Ti0>0 Li0>1 Li1>7 To0<0 Ro0<15 ]
  led g38 (.I(w24));   //: @(780,393) /sn:0 /R:2 /w:[ 7 ] /type:2
  //: dip g27 (w12) @(920,153) /sn:0 /w:[ 0 ] /st:0
  //: joint g37 (w11) @(843, 184) /w:[ 2 -1 4 1 ]
  mux g13 (.I0(w24), .I1(w25), .S(w14), .Z(w22));   //: @(817,271) /sn:0 /R:1 /w:[ 5 3 1 0 ] /ss:1 /do:1

endmodule

module Read(SignExOut, SignExIn, RegDst, R1, R2, WR, RD2, WriteData, RD1, clk, clr, RegWrite);
//: interface  /sz:(162, 244) /bd:[ Ti0>RegWrite(85/162) Ti1>RegWrite(85/162) Ti2>RegWrite(85/162) Li0>R1[4:0](34/244) Li1>R2[4:0](65/244) Li2>WR[4:0](97/244) Li3>RegDst(122/244) Li4>WriteData[31:0](153/244) Li5>SignExIn[15:0](200/244) Li6>SignExIn[15:0](200/244) Li7>WriteData[31:0](153/244) Li8>RegDst(122/244) Li9>WR[4:0](97/244) Li10>R2[4:0](65/244) Li11>R1[4:0](34/244) Li12>SignExIn[15:0](200/244) Li13>WriteData[31:0](153/244) Li14>RegDst(122/244) Li15>WR[4:0](97/244) Li16>R2[4:0](65/244) Li17>R1[4:0](34/244) Bi0>clk(55/162) Bi1>clr(111/162) Bi2>clr(111/162) Bi3>clk(55/162) Bi4>clr(111/162) Bi5>clk(55/162) Ro0<RD1[31:0](49/244) Ro1<RD2[31:0](126/244) Ro2<SignExOut[31:0](205/244) Ro3<SignExOut[31:0](205/244) Ro4<RD2[31:0](126/244) Ro5<RD1[31:0](49/244) Ro6<SignExOut[31:0](205/244) Ro7<RD2[31:0](126/244) Ro8<RD1[31:0](49/244) ]
input [4:0] WR;    //: /sn:0 {0}(411,219)(464,219){1}
input [31:0] WriteData;    //: /sn:0 {0}(500,249)(532,249){1}
input [4:0] R2;    //: /sn:0 {0}(412,173)(435,173){1}
//: {2}(439,173)(532,173){3}
//: {4}(437,175)(437,199)(464,199){5}
output [31:0] SignExOut;    //: /sn:0 {0}(718,440)(637,440){1}
output [31:0] RD2;    //: /sn:0 {0}(720,240)(681,240){1}
input [4:0] R1;    //: /sn:0 {0}(411,133)(532,133){1}
input RegDst;    //: /sn:0 {0}(463,271)(480,271)(480,232){1}
input clr;    //: /sn:0 {0}(585,65)(599,65)(599,100){1}
input RegWrite;    //: /sn:0 {0}(565,324)(573,324)(573,284){1}
input clk;    //: /sn:0 {0}(624,322)(641,322)(641,284){1}
output [31:0] RD1;    //: /sn:0 {0}(724,148)(681,148){1}
input [15:0] SignExIn;    //: /sn:0 {0}(499,441)(571,441){1}
wire [4:0] w12;    //: /sn:0 /dp:1 {0}(493,209)(532,209){1}
//: enddecls

  //: output g4 (SignExOut) @(715,440) /sn:0 /w:[ 0 ]
  //: joint g8 (R2) @(437, 173) /w:[ 2 -1 1 4 ]
  //: input g3 (SignExIn) @(497,441) /sn:0 /w:[ 0 ]
  mux g2 (.I0(WR), .I1(R2), .S(RegDst), .Z(w12));   //: @(480,209) /sn:0 /R:1 /w:[ 1 5 1 0 ] /ss:0 /do:0
  Sign_extend g1 (.in(SignExIn), .out(SignExOut));   //: @(572, 404) /sz:(64, 66) /sn:0 /p:[ Li0>1 Ro0<1 ]
  //: input g10 (RegDst) @(461,271) /sn:0 /w:[ 0 ]
  //: input g6 (R1) @(409,133) /sn:0 /w:[ 0 ]
  //: input g7 (R2) @(410,173) /sn:0 /w:[ 0 ]
  //: input g9 (WR) @(409,219) /sn:0 /w:[ 0 ]
  //: output g12 (RD2) @(717,240) /sn:0 /w:[ 0 ]
  //: input g5 (WriteData) @(498,249) /sn:0 /w:[ 0 ]
  //: output g11 (RD1) @(721,148) /sn:0 /w:[ 0 ]
  //: input g14 (clk) @(622,322) /sn:0 /w:[ 0 ]
  BRegs32x32 g0 (.clr(clr), .Read1(R1), .Read2(R2), .Write(w12), .WriteData(WriteData), .clk(clk), .RegWrite(RegWrite), .Data1(RD1), .Data2(RD2));   //: @(533, 101) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>1 Li1>3 Li2>1 Li3>1 Bi0>1 Bi1>1 Ro0<1 Ro1<1 ]
  //: input g15 (clr) @(583,65) /sn:0 /w:[ 0 ]
  //: input g13 (RegWrite) @(563,324) /sn:0 /w:[ 0 ]

endmodule

module Sign_extend(out, in);
//: interface  /sz:(64, 66) /bd:[ Li0>in[15:0](37/66) Ro0<out[31:0](36/66) ]
input [15:0] in;    //: /sn:0 {0}(441,165)(464,165)(464,166){1}
//: {2}(464,167)(464,350){3}
//: {4}(464,351)(464,359){5}
output [31:0] out;    //: /sn:0 {0}(606,266)(571,266){1}
wire [14:0] w0;    //: /sn:0 {0}(468,351)(565,351){1}
wire w18;    //: /sn:0 {0}(565,181)(473,181){1}
//: {2}(471,179)(471,167)(468,167){3}
//: {4}(471,183)(471,199){5}
//: {6}(473,201)(521,201){7}
//: {8}(525,201)(565,201){9}
//: {10}(523,199)(523,191)(565,191){11}
//: {12}(471,203)(471,219){13}
//: {14}(473,221)(521,221){15}
//: {16}(525,221)(565,221){17}
//: {18}(523,219)(523,211)(565,211){19}
//: {20}(471,223)(471,239){21}
//: {22}(473,241)(521,241){23}
//: {24}(525,241)(565,241){25}
//: {26}(523,239)(523,231)(565,231){27}
//: {28}(471,243)(471,259){29}
//: {30}(473,261)(521,261){31}
//: {32}(525,261)(565,261){33}
//: {34}(523,259)(523,251)(565,251){35}
//: {36}(471,263)(471,279){37}
//: {38}(473,281)(520,281){39}
//: {40}(524,281)(565,281){41}
//: {42}(522,279)(522,271)(565,271){43}
//: {44}(471,283)(471,299){45}
//: {46}(473,301)(520,301){47}
//: {48}(524,301)(565,301){49}
//: {50}(522,299)(522,291)(565,291){51}
//: {52}(471,303)(471,319){53}
//: {54}(473,321)(519,321){55}
//: {56}(523,321)(565,321){57}
//: {58}(521,319)(521,311)(565,311){59}
//: {60}(471,323)(471,339){61}
//: {62}(473,341)(519,341){63}
//: {64}(523,341)(565,341){65}
//: {66}(521,339)(521,331)(565,331){67}
//: {68}(471,343)(471,348){69}
//: enddecls

  tran g4(.Z(w18), .I(in[15]));   //: @(462,167) /sn:0 /R:2 /w:[ 3 2 1 ] /ss:1
  //: joint g8 (w18) @(521, 321) /w:[ 56 58 55 -1 ]
  tran g3(.Z(w0), .I(in[14:0]));   //: @(462,351) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: joint g16 (w18) @(523, 241) /w:[ 24 26 23 -1 ]
  //: joint g17 (w18) @(471, 221) /w:[ 14 13 -1 20 ]
  concat g2 (.I0(w0), .I1(w18), .I2(w18), .I3(w18), .I4(w18), .I5(w18), .I6(w18), .I7(w18), .I8(w18), .I9(w18), .I10(w18), .I11(w18), .I12(w18), .I13(w18), .I14(w18), .I15(w18), .I16(w18), .I17(w18), .Z(out));   //: @(570,266) /sn:0 /w:[ 1 65 67 57 59 49 51 41 43 33 35 25 27 17 19 9 11 0 1 ] /dr:0
  //: output g1 (out) @(603,266) /sn:0 /w:[ 0 ]
  //: joint g18 (w18) @(523, 221) /w:[ 16 18 15 -1 ]
  //: joint g10 (w18) @(522, 301) /w:[ 48 50 47 -1 ]
  //: joint g6 (w18) @(521, 341) /w:[ 64 66 63 -1 ]
  //: joint g7 (w18) @(471, 321) /w:[ 54 53 -1 60 ]
  //: joint g9 (w18) @(471, 301) /w:[ 46 45 -1 52 ]
  //: joint g12 (w18) @(522, 281) /w:[ 40 42 39 -1 ]
  //: joint g5 (w18) @(471, 341) /w:[ 62 61 -1 68 ]
  //: joint g11 (w18) @(471, 281) /w:[ 38 37 -1 44 ]
  //: joint g14 (w18) @(523, 261) /w:[ 32 34 31 -1 ]
  //: joint g19 (w18) @(471, 201) /w:[ 6 5 -1 12 ]
  //: joint g21 (w18) @(471, 181) /w:[ 1 2 -1 4 ]
  //: joint g20 (w18) @(523, 201) /w:[ 8 10 7 -1 ]
  //: input g0 (in) @(439,165) /sn:0 /w:[ 0 ]
  //: joint g15 (w18) @(471, 241) /w:[ 22 21 -1 28 ]
  //: joint g13 (w18) @(471, 261) /w:[ 30 29 -1 36 ]

endmodule
