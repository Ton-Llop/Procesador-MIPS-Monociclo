//: version "1.8.7"

module ALU(B, AluResult, AluOp, Z, A);
//: interface  /sz:(40, 40) /bd:[ ]
input [31:0] B;    //: /sn:0 {0}(238,220)(301,220)(301,308){1}
//: {2}(303,310)(390,310)(390,367)(405,367){3}
//: {4}(301,312)(301,345)(307,345)(307,367)(313,367){5}
supply0 [30:0] w4;    //: /sn:0 {0}(520,272)(520,298)(528,298)(528,315)(539,315){1}
input [31:0] A;    //: /sn:0 /dp:1 {0}(427,167)(411,167)(411,153)(408,153){1}
//: {2}(404,153)(365,153){3}
//: {4}(361,153)(239,153){5}
//: {6}(363,155)(363,242)(476,242){7}
//: {8}(406,155)(406,200)(445,200){9}
output Z;    //: /sn:0 {0}(764,218)(754,218)(754,217)(715,217){1}
output [31:0] AluResult;    //: /sn:0 {0}(736,286)(672,286)(672,254){1}
//: {2}(672,250)(672,217)(694,217){3}
//: {4}(670,252)(629,252){5}
input [3:0] AluOp;    //: /sn:0 {0}(231,446)(394,446){1}
//: {2}(395,446)(469,446)(469,447)(543,447){3}
//: {4}(544,447)(646,447){5}
wire [31:0] w13;    //: /sn:0 /dp:1 {0}(600,270)(564,270)(564,320)(545,320){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(427,172)(422,172)(422,265)(442,265)(442,280){1}
//: {2}(440,282)(436,282)(436,195)(445,195){3}
//: {4}(442,284)(442,347)(456,347)(456,355){5}
//: {6}(458,357)(470,357)(470,274)(476,274){7}
//: {8}(454,357)(434,357){9}
wire [31:0] w12;    //: /sn:0 /dp:3 {0}(600,258)(511,258){1}
//: {2}(510,258)(505,258){3}
wire w1;    //: /sn:0 {0}(511,262)(511,325)(539,325){1}
wire [31:0] po;    //: /sn:0 {0}(405,347)(374,347)(374,367)(329,367){1}
wire [31:0] w17;    //: /sn:0 /dp:1 {0}(466,197)(562,197)(562,246)(600,246){1}
wire [1:0] w14;    //: /sn:0 /dp:1 {0}(544,442)(544,361)(616,361)(616,275){1}
wire w2;    //: /sn:0 {0}(421,380)(421,393){1}
//: {2}(423,395)(446,395)(446,224)(490,224)(490,234){3}
//: {4}(421,397)(421,434)(395,434)(395,441){5}
wire [31:0] w15;    //: /sn:0 /dp:1 {0}(448,169)(594,169)(594,234)(600,234){1}
wire w5;    //: /sn:0 /dp:1 {0}(490,337)(490,282){1}
//: enddecls

  not g4 (.I(B), .Z(po));   //: @(319,367) /sn:0 /w:[ 5 1 ]
  mux g8 (.I0(w15), .I1(w17), .I2(w12), .I3(w13), .S(w14), .Z(AluResult));   //: @(616,252) /sn:0 /R:1 /w:[ 1 1 0 0 1 5 ] /ss:0 /do:1
  mux g3 (.I0(B), .I1(po), .S(w2), .Z(w3));   //: @(421,357) /sn:0 /R:1 /w:[ 3 0 0 9 ] /ss:0 /do:0
  //: joint g16 (w2) @(421, 395) /w:[ 2 1 -1 4 ]
  concat g17 (.I0(w1), .I1(w4), .Z(w13));   //: @(544,320) /sn:0 /w:[ 1 1 1 ] /dr:0
  //: joint g2 (B) @(301, 310) /w:[ 2 1 -1 4 ]
  nor g23 (.I0(AluResult), .Z(Z));   //: @(705,217) /sn:0 /w:[ 3 1 ]
  //: input g1 (B) @(236,220) /sn:0 /w:[ 0 ]
  //: output g24 (AluResult) @(733,286) /sn:0 /w:[ 0 ]
  tran g18(.Z(w1), .I(w12[31]));   //: @(511,256) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  and g10 (.I0(A), .I1(w3), .Z(w15));   //: @(438,169) /sn:0 /w:[ 0 0 0 ]
  add g6 (.A(w3), .B(A), .S(w12), .CI(w2), .CO(w5));   //: @(492,258) /sn:0 /R:1 /w:[ 7 7 3 3 1 ]
  tran g9(.Z(w2), .I(AluOp[2]));   //: @(395,444) /sn:0 /R:1 /w:[ 5 1 2 ] /ss:0
  tran g7(.Z(w14), .I(AluOp[1:0]));   //: @(544,445) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:0
  //: joint g22 (AluResult) @(672, 252) /w:[ -1 2 4 1 ]
  //: joint g12 (w3) @(442, 282) /w:[ -1 1 2 4 ]
  //: input g5 (AluOp) @(229,446) /sn:0 /w:[ 0 ]
  or g11 (.I0(w3), .I1(A), .Z(w17));   //: @(456,197) /sn:0 /w:[ 3 9 0 ]
  //: joint g14 (w3) @(456, 357) /w:[ 6 5 8 -1 ]
  //: supply0 g19 (w4) @(520,266) /sn:0 /R:2 /w:[ 0 ]
  //: output g21 (Z) @(761,218) /sn:0 /w:[ 0 ]
  led g20 (.I(w5));   //: @(490,344) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: input g0 (A) @(237,153) /sn:0 /w:[ 5 ]
  //: joint g15 (A) @(363, 153) /w:[ 3 -1 4 6 ]
  //: joint g13 (A) @(406, 153) /w:[ 1 -1 2 8 ]

endmodule

module main;    //: root_module
wire [3:0] w7;    //: /sn:0 /dp:1 {0}(916,235)(916,262){1}
wire w4;    //: /sn:0 {0}(1043,250)(1043,316)(995,316){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(601,251)(601,290)(822,290){1}
wire w10;    //: /sn:0 {0}(23354,-6430)(23354,-6420){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(488,307)(488,316)(822,316){1}
wire w8;    //: /sn:0 {0}(23302,-6422)(23302,-6412){1}
wire w2;    //: /sn:0 {0}(23290,-6401)(23290,-6391){1}
wire [31:0] w5;    //: /sn:0 {0}(1136,331)(1136,355)(995,355){1}
//: enddecls

  led g4 (.I(w5));   //: @(1136,324) /sn:0 /w:[ 0 ] /type:2
  ALU g3 (.AluOp(w7), .B(w1), .A(w0), .AluResult(w5), .Z(w4));   //: @(823, 263) /sz:(171, 157) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<1 Ro1<1 ]
  //: dip g1 (w1) @(488,297) /sn:0 /w:[ 0 ] /st:5
  //: switch g10 (w2) @(23290,-6414) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: dip g6 (w7) @(916,225) /sn:0 /w:[ 0 ] /st:0
  //: switch g12 (w10) @(23354,-6443) /sn:0 /R:3 /w:[ 0 ] /st:0
  led g5 (.I(w4));   //: @(1043,243) /sn:0 /w:[ 0 ] /type:0
  //: switch g11 (w8) @(23302,-6435) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: dip g0 (w0) @(601,241) /sn:0 /w:[ 0 ] /st:5

endmodule
