//: version "1.8.7"

module memoria(RD, WD, Addr, MemRead, MemWrite, clk);
//: interface  /sz:(297, 200) /bd:[ Ti0>MemWrite(147/297) Li0>WD[31:0](133/200) Li1>Addr[31:0](37/200) Bi0>clk(224/297) Bi1>MemRead(133/297) Ro0<RD[31:0](82/200) ]
supply0 w0;    //: /sn:0 {0}(715,297)(715,278){1}
input [31:0] Addr;    //: /sn:0 {0}(668,253)(704,253){1}
input [31:0] WD;    //: /sn:0 /dp:1 {0}(786,224)(786,201)(771,201){1}
input MemWrite;    //: /sn:0 {0}(623,163)(718,163){1}
//: {2}(722,163)(809,163)(809,232)(791,232){3}
//: {4}(720,165)(720,181){5}
input clk;    //: /sn:0 {0}(637,147)(725,147)(725,181){1}
output [31:0] RD;    //: /sn:0 {0}(833,251)(788,251){1}
//: {2}(786,249)(786,240){3}
//: {4}(784,251)(739,251){5}
input MemRead;    //: /sn:0 {0}(683,339)(729,339)(729,278){1}
wire w9;    //: /sn:0 {0}(722,202)(722,228){1}
//: enddecls

  //: output g4 (RD) @(830,251) /sn:0 /w:[ 0 ]
  bufif1 g8 (.Z(RD), .I(WD), .E(MemWrite));   //: @(786,230) /sn:0 /R:3 /w:[ 3 0 3 ]
  //: input g3 (WD) @(769,201) /sn:0 /w:[ 1 ]
  //: supply0 g2 (w0) @(715,303) /sn:0 /w:[ 0 ]
  //: input g1 (Addr) @(666,253) /sn:0 /w:[ 0 ]
  //: joint g10 (MemWrite) @(720, 163) /w:[ 2 -1 1 4 ]
  //: input g6 (MemRead) @(681,339) /sn:0 /w:[ 0 ]
  //: input g7 (MemWrite) @(621,163) /sn:0 /w:[ 0 ]
  nand g9 (.I0(clk), .I1(MemWrite), .Z(w9));   //: @(722,192) /sn:0 /R:3 /w:[ 1 5 0 ]
  //: input g5 (clk) @(635,147) /sn:0 /w:[ 0 ]
  //: joint g11 (RD) @(786, 251) /w:[ 1 2 4 -1 ]
  ram g0 (.A(Addr), .D(RD), .WE(w9), .OE(!MemRead), .CS(w0));   //: @(722,252) /sn:0 /w:[ 1 5 1 1 1 ]

endmodule

module main;    //: root_module
wire [31:0] w4;    //: /sn:0 {0}(476,330)(476,350)(530,350){1}
wire [31:0] w3;    //: /sn:0 {0}(469,244)(469,254)(530,254){1}
wire w0;    //: /sn:0 {0}(653,171)(678,171)(678,216){1}
wire w1;    //: /sn:0 {0}(638,455)(664,455)(664,418){1}
wire w2;    //: /sn:0 {0}(752,458)(755,458)(755,418){1}
wire [31:0] w5;    //: /sn:0 {0}(919,290)(919,299)(829,299){1}
//: enddecls

  //: dip g4 (w3) @(469,234) /sn:0 /w:[ 0 ] /st:0
  //: switch g3 (w2) @(735,458) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w1) @(621,455) /sn:0 /w:[ 0 ] /st:1
  //: switch g1 (w0) @(636,171) /sn:0 /w:[ 0 ] /st:0
  led g6 (.I(w5));   //: @(919,283) /sn:0 /w:[ 0 ] /type:2
  //: dip g5 (w4) @(476,320) /sn:0 /w:[ 0 ] /st:5397
  memoria g0 (.MemWrite(w0), .WD(w4), .Addr(w3), .clk(w2), .MemRead(w1), .RD(w5));   //: @(531, 217) /sz:(297, 200) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bi0>1 Bi1>1 Ro0<1 ]

endmodule
