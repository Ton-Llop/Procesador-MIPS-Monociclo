//: version "1.8.7"

module jump(SignXtended, dir, PCNext, jump, PCSrc, inm26);
//: interface  /sz:(121, 80) /bd:[ Ti0>jump(74/121) Li0>PCNext[31:0](51/80) Li1>inm26[25:0](19/80) Bi0>PCSrc(85/121) Bi1>SignXtended[31:0](37/121) Ro0<dir[31:0](36/80) ]
input jump;    //: /sn:0 {0}(503,158)(503,124){1}
input PCSrc;    //: /sn:0 /dp:1 {0}(433,134)(433,180){1}
input [25:0] inm26;    //: /sn:0 {0}(139,76)(272,76){1}
supply0 w3;    //: /sn:0 {0}(328,47)(328,97){1}
output [31:0] dir;    //: /sn:0 /dp:1 {0}(516,101)(568,101){1}
input [31:0] PCNext;    //: /sn:0 /dp:1 {0}(417,101)(353,101)(353,83)(301,83)(301,103){1}
//: {2}(303,105)(314,105){3}
//: {4}(299,105)(203,105){5}
//: {6}(202,105)(139,105){7}
input [31:0] SignXtended;    //: /sn:0 /dp:1 {0}(314,137)(292,137)(292,175){1}
wire w6;    //: /sn:0 /dp:1 {0}(328,145)(328,155){1}
wire [31:0] w7;    //: /sn:0 {0}(417,121)(343,121){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(487,111)(446,111){1}
wire [5:0] w1;    //: /sn:0 {0}(203,100)(203,66)(272,66){1}
wire [31:0] w2;    //: /sn:0 {0}(278,71)(461,71)(461,91)(487,91){1}
//: enddecls

  concat g4 (.I0(inm26), .I1(w1), .Z(w2));   //: @(277,71) /sn:0 /w:[ 1 1 0 ] /dr:0
  mux g8 (.I0(PCNext), .I1(w7), .S(PCSrc), .Z(w0));   //: @(433,111) /sn:0 /R:1 /w:[ 0 0 0 1 ] /ss:0 /do:1
  //: input g3 (SignXtended) @(292,177) /sn:0 /R:1 /w:[ 1 ]
  //: output g2 (dir) @(565,101) /sn:0 /w:[ 1 ]
  //: input g1 (PCNext) @(137,105) /sn:0 /w:[ 7 ]
  //: joint g10 (PCNext) @(301, 105) /w:[ 2 1 4 -1 ]
  add g6 (.A(SignXtended), .B(PCNext), .S(w7), .CI(w3), .CO(w6));   //: @(330,121) /sn:0 /R:1 /w:[ 0 3 1 1 0 ]
  mux g7 (.I0(w0), .I1(w2), .S(jump), .Z(dir));   //: @(503,101) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:0 /do:0
  //: input g9 (jump) @(503,160) /sn:0 /R:1 /w:[ 0 ]
  //: supply0 g12 (w3) @(328,41) /sn:0 /R:2 /w:[ 0 ]
  tran g5(.Z(w1), .I(PCNext[31:26]));   //: @(203,103) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:0
  //: input g11 (PCSrc) @(433,182) /sn:0 /R:1 /w:[ 1 ]
  //: input g0 (inm26) @(137,76) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [31:0] w6;    //: /sn:0 {0}(187,182)(187,196)(339,196){1}
wire [15:0] w7;    //: /sn:0 {0}(215,276)(215,293)(271,293){1}
wire [31:0] w4;    //: /sn:0 {0}(576,172)(576,181)(462,181){1}
wire w3;    //: /sn:0 {0}(422,264)(425,264)(425,226){1}
wire [31:0] w1;    //: /sn:0 {0}(337,292)(377,292)(377,226){1}
wire w2;    //: /sn:0 {0}(405,110)(414,110)(414,144){1}
wire [25:0] w5;    //: /sn:0 {0}(248,145)(248,164)(339,164){1}
//: enddecls

  led g4 (.I(w4));   //: @(576,165) /sn:0 /w:[ 0 ] /type:2
  //: switch g3 (w3) @(405,264) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w2) @(388,110) /sn:0 /w:[ 0 ] /st:0
  Sign_extend g1 (.in(w7), .out(w1));   //: @(272, 256) /sz:(64, 66) /sn:0 /p:[ Li0>1 Ro0<0 ]
  //: dip g6 (w6) @(187,172) /sn:0 /w:[ 0 ] /st:-52428800
  //: dip g7 (w7) @(215,266) /sn:0 /w:[ 0 ] /st:4369
  //: dip g5 (w5) @(248,135) /sn:0 /w:[ 0 ] /st:4194303
  jump g0 (.jump(w2), .PCNext(w6), .inm26(w5), .PCSrc(w3), .SignXtended(w1), .dir(w4));   //: @(340, 145) /sz:(121, 80) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bi0>1 Bi1>1 Ro0<1 ]

endmodule

module Sign_extend(out, in);
//: interface  /sz:(64, 66) /bd:[ Li0>in[15:0](37/66) Ro0<out[31:0](36/66) ]
input [15:0] in;    //: /sn:0 {0}(441,165)(464,165)(464,166){1}
//: {2}(464,167)(464,350){3}
//: {4}(464,351)(464,359){5}
output [31:0] out;    //: /sn:0 {0}(606,266)(571,266){1}
wire [14:0] w0;    //: /sn:0 {0}(468,351)(565,351){1}
wire w18;    //: /sn:0 {0}(565,181)(473,181){1}
//: {2}(471,179)(471,167)(468,167){3}
//: {4}(471,183)(471,199){5}
//: {6}(473,201)(521,201){7}
//: {8}(525,201)(565,201){9}
//: {10}(523,199)(523,191)(565,191){11}
//: {12}(471,203)(471,219){13}
//: {14}(473,221)(521,221){15}
//: {16}(525,221)(565,221){17}
//: {18}(523,219)(523,211)(565,211){19}
//: {20}(471,223)(471,239){21}
//: {22}(473,241)(521,241){23}
//: {24}(525,241)(565,241){25}
//: {26}(523,239)(523,231)(565,231){27}
//: {28}(471,243)(471,259){29}
//: {30}(473,261)(521,261){31}
//: {32}(525,261)(565,261){33}
//: {34}(523,259)(523,251)(565,251){35}
//: {36}(471,263)(471,279){37}
//: {38}(473,281)(520,281){39}
//: {40}(524,281)(565,281){41}
//: {42}(522,279)(522,271)(565,271){43}
//: {44}(471,283)(471,299){45}
//: {46}(473,301)(520,301){47}
//: {48}(524,301)(565,301){49}
//: {50}(522,299)(522,291)(565,291){51}
//: {52}(471,303)(471,319){53}
//: {54}(473,321)(519,321){55}
//: {56}(523,321)(565,321){57}
//: {58}(521,319)(521,311)(565,311){59}
//: {60}(471,323)(471,339){61}
//: {62}(473,341)(519,341){63}
//: {64}(523,341)(565,341){65}
//: {66}(521,339)(521,331)(565,331){67}
//: {68}(471,343)(471,348){69}
//: enddecls

  tran g4(.Z(w18), .I(in[15]));   //: @(462,167) /sn:0 /R:2 /w:[ 3 2 1 ] /ss:1
  //: joint g8 (w18) @(521, 321) /w:[ 56 58 55 -1 ]
  tran g3(.Z(w0), .I(in[14:0]));   //: @(462,351) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: joint g16 (w18) @(523, 241) /w:[ 24 26 23 -1 ]
  //: joint g17 (w18) @(471, 221) /w:[ 14 13 -1 20 ]
  concat g2 (.I0(w0), .I1(w18), .I2(w18), .I3(w18), .I4(w18), .I5(w18), .I6(w18), .I7(w18), .I8(w18), .I9(w18), .I10(w18), .I11(w18), .I12(w18), .I13(w18), .I14(w18), .I15(w18), .I16(w18), .I17(w18), .Z(out));   //: @(570,266) /sn:0 /w:[ 1 65 67 57 59 49 51 41 43 33 35 25 27 17 19 9 11 0 1 ] /dr:0
  //: output g1 (out) @(603,266) /sn:0 /w:[ 0 ]
  //: joint g18 (w18) @(523, 221) /w:[ 16 18 15 -1 ]
  //: joint g10 (w18) @(522, 301) /w:[ 48 50 47 -1 ]
  //: joint g6 (w18) @(521, 341) /w:[ 64 66 63 -1 ]
  //: joint g7 (w18) @(471, 321) /w:[ 54 53 -1 60 ]
  //: joint g9 (w18) @(471, 301) /w:[ 46 45 -1 52 ]
  //: joint g12 (w18) @(522, 281) /w:[ 40 42 39 -1 ]
  //: joint g5 (w18) @(471, 341) /w:[ 62 61 -1 68 ]
  //: joint g11 (w18) @(471, 281) /w:[ 38 37 -1 44 ]
  //: joint g14 (w18) @(523, 261) /w:[ 32 34 31 -1 ]
  //: joint g19 (w18) @(471, 201) /w:[ 6 5 -1 12 ]
  //: joint g21 (w18) @(471, 181) /w:[ 1 2 -1 4 ]
  //: joint g20 (w18) @(523, 201) /w:[ 8 10 7 -1 ]
  //: input g0 (in) @(439,165) /sn:0 /w:[ 0 ]
  //: joint g15 (w18) @(471, 241) /w:[ 22 21 -1 28 ]
  //: joint g13 (w18) @(471, 261) /w:[ 30 29 -1 36 ]

endmodule
