//: version "1.8.7"

module Fetch(Inst, Reset, Clk, PCIn, PCOut);
//: interface  /sz:(107, 96) /bd:[ Ti0>PCIn[31:0](76/107) Li0>Clk(65/96) Li1>Reset(22/96) To0<PCOut[31:0](28/107) Ro0<Inst[31:0](49/96) ]
supply0 w13;    //: /sn:0 {0}(348,222)(348,195){1}
output [31:0] PCOut;    //: /sn:0 /dp:1 {0}(429,76)(482,76){1}
input Clk;    //: /sn:0 {0}(188,208)(238,208)(238,185){1}
output [31:0] Inst;    //: /sn:0 {0}(427,168)(365,168){1}
input [31:0] PCIn;    //: /sn:0 {0}(148,147)(227,147){1}
input Reset;    //: /sn:0 {0}(182,91)(233,91)(233,109){1}
supply0 w14;    //: /sn:0 {0}(258,73)(258,99)(243,99)(243,109){1}
supply0 w15;    //: /sn:0 {0}(439,39)(414,39)(414,52){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(352,46)(352,60)(400,60){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(248,147)(301,147){1}
//: {2}(305,147)(326,147)(326,170)(330,170){3}
//: {4}(303,145)(303,92)(400,92){5}
wire w12;    //: /sn:0 {0}(414,100)(414,110){1}
//: enddecls

  //: output g8 (Inst) @(424,168) /sn:0 /w:[ 0 ]
  //: supply0 g4 (w14) @(258,67) /sn:0 /R:2 /w:[ 0 ]
  //: supply0 g3 (w13) @(348,228) /sn:0 /w:[ 0 ]
  add g2 (.A(w3), .B(w0), .S(PCOut), .CI(w15), .CO(w12));   //: @(416,76) /sn:0 /R:1 /w:[ 5 1 0 1 0 ]
  register g1 (.Q(w3), .D(PCIn), .EN(w14), .CLR(!Reset), .CK(Clk));   //: @(238,147) /sn:0 /R:1 /w:[ 0 1 1 1 1 ]
  //: input g10 (Reset) @(180,91) /sn:0 /w:[ 0 ]
  //: joint g6 (w3) @(303, 147) /w:[ 2 4 1 -1 ]
  //: input g9 (Clk) @(186,208) /sn:0 /w:[ 0 ]
  //: dip g7 (w0) @(352,36) /sn:0 /w:[ 0 ] /st:1
  //: input g12 (PCIn) @(146,147) /sn:0 /w:[ 0 ]
  //: supply0 g5 (w15) @(445,39) /sn:0 /R:1 /w:[ 0 ]
  //: output g11 (PCOut) @(479,76) /sn:0 /w:[ 1 ]
  rom g0 (.A(w3), .D(Inst), .OE(w13));   //: @(348,169) /sn:0 /w:[ 3 1 1 ]

endmodule

module main;    //: root_module
wire w13;    //: /sn:0 {0}(145,240)(220,240)(220,139)(230,139){1}
wire w0;    //: /sn:0 {0}(171,96)(230,96){1}
wire [31:0] w1;    //: /sn:0 {0}(440,109)(440,123)(339,123){1}
wire [31:0] PCIn;    //: /sn:0 {0}(307,73)(307,45)(259,45)(259,73){1}
//: enddecls

  clock g3 (.Z(w13));   //: @(132,240) /sn:0 /w:[ 0 ] /omega:2000 /phi:0 /duty:50
  led g1 (.I(w1));   //: @(440,102) /sn:0 /w:[ 0 ] /type:2
  Fetch g12 (.PCIn(PCIn), .Clk(w13), .Reset(w0), .PCOut(PCIn), .Inst(w1));   //: @(231, 74) /sz:(107, 96) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 To0<1 Ro0<1 ]
  //: switch g0 (w0) @(154,96) /sn:0 /w:[ 0 ] /st:0

endmodule
