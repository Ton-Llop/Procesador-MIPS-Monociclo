//: version "1.8.7"

module jump(SignXtended, dir, PCNext, jump, PCSrc, inm26);
//: interface  /sz:(121, 80) /bd:[ Ti0>jump(74/121) Li0>PCNext[31:0](51/80) Li1>inm26[25:0](19/80) Bi0>PCSrc(85/121) Bi1>SignXtended[31:0](37/121) Ro0<dir[31:0](36/80) ]
input jump;    //: /sn:0 {0}(503,158)(503,124){1}
input PCSrc;    //: /sn:0 /dp:1 {0}(433,134)(433,124)(448,124)(448,180){1}
input [25:0] inm26;    //: /sn:0 {0}(139,76)(272,76){1}
supply0 w3;    //: /sn:0 {0}(328,47)(328,57)(343,57)(353,47)(353,62)(343,102)(328,102)(328,112){1}
output [31:0] dir;    //: /sn:0 /dp:1 {0}(516,101)(568,101){1}
input [31:0] PCNext;    //: /sn:0 /dp:1 {0}(417,101)(353,101)(353,83)(301,83)(301,103){1}
//: {2}(303,105)(314,105){3}
//: {4}(299,105)(203,105){5}
//: {6}(202,105)(139,105){7}
input [31:0] SignXtended;    //: /sn:0 /dp:1 {0}(314,137)(292,137)(292,175){1}
wire w6;    //: /sn:0 /dp:1 {0}(328,145)(328,155){1}
wire [31:0] w7;    //: /sn:0 {0}(417,121)(343,121){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(487,111)(446,111){1}
wire [5:0] w1;    //: /sn:0 {0}(203,99)(203,66)(272,66){1}
wire [31:0] w2;    //: /sn:0 {0}(278,71)(461,71)(461,91)(487,91){1}
//: enddecls

  concat g4 (.I0(inm26), .I1(w1), .Z(w2));   //: @(277,71) /sn:0 /w:[ 1 1 0 ] /dr:0
  mux g8 (.I0(PCNext), .I1(w7), .S(PCSrc), .Z(w0));   //: @(433,111) /sn:0 /R:1 /w:[ 0 0 0 1 ] /ss:1 /do:1
  //: input g3 (SignXtended) @(292,177) /sn:0 /R:1 /w:[ 1 ]
  //: output g2 (dir) @(565,101) /sn:0 /w:[ 1 ]
  //: input g1 (PCNext) @(137,105) /sn:0 /w:[ 7 ]
  //: joint g10 (PCNext) @(301, 105) /w:[ 2 1 4 -1 ]
  add g6 (.A(SignXtended), .B(PCNext), .S(w7), .CI(w3), .CO(w6));   //: @(330,121) /sn:0 /R:1 /w:[ 0 3 1 1 0 ]
  mux g7 (.I0(w0), .I1(w2), .S(jump), .Z(dir));   //: @(503,101) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:1 /do:1
  //: input g9 (jump) @(503,160) /sn:0 /R:1 /w:[ 0 ]
  //: supply0 g12 (w3) @(328,41) /sn:0 /R:2 /w:[ 0 ]
  //: input g11 (PCSrc) @(433,182) /sn:0 /R:1 /w:[ 1 ]
  tran g5(.Z(w1), .I(PCNext[31:26]));   //: @(203,103) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:0
  //: input g0 (inm26) @(137,76) /sn:0 /w:[ 0 ]

endmodule

module UC(Jump, MemWrite, RegWrite, MemRead, ALUCtrl, ALUSrc, MemToReg, Branch, Ins, RegDst);
//: interface  /sz:(132, 331) /bd:[ Li0>Ins[31:0](151/331) Ro0<RegDst(36/331) Ro1<Branch(70/331) Ro2<Jump(107/331) Ro3<MemRead(138/331) Ro4<MemToReg(171/331) Ro5<ALUCtrl[3:0](203/331) Ro6<MemWrite(232/331) Ro7<ALUSrc(259/331) Ro8<RegWrite(288/331) ]
output Branch;    //: /sn:0 /dp:1 {0}(378,101)(378,263)(512,263){1}
//: {2}(514,261)(514,254)(535,254){3}
//: {4}(514,265)(514,273){5}
output [3:0] ALUCtrl;    //: /sn:0 /dp:1 {0}(414,51)(434,51){1}
output MemWrite;    //: /sn:0 /dp:1 {0}(463,274)(463,271){1}
//: {2}(465,269)(473,269)(473,153)(556,153){3}
//: {4}(560,153)(725,153){5}
//: {6}(558,155)(558,189)(658,189){7}
//: {8}(463,267)(463,252){9}
output ALUSrc;    //: /sn:0 /dp:1 {0}(679,187)(715,187)(715,185)(726,185){1}
input [31:0] Ins;    //: /sn:0 {0}(202,330)(213,330){1}
//: {2}(217,330)(250,330)(250,335){3}
//: {4}(250,336)(250,344){5}
//: {6}(250,345)(250,352){7}
//: {8}(250,353)(250,360){9}
//: {10}(250,361)(250,368){11}
//: {12}(250,369)(250,376){13}
//: {14}(250,377)(250,487){15}
//: {16}(215,328)(215,187){17}
//: {18}(215,186)(215,164){19}
//: {20}(215,163)(215,128){21}
//: {22}(215,127)(215,107){23}
//: {24}(215,106)(215,65){25}
output RegDst;    //: /sn:0 /dp:1 {0}(334,109)(334,266)(353,266){1}
//: {2}(357,266)(363,266)(363,275){3}
//: {4}(355,264)(355,256)(354,256)(354,246){5}
//: {6}(356,244)(366,244)(366,243)(373,243){7}
//: {8}(354,242)(354,225){9}
//: {10}(356,223)(659,223){11}
//: {12}(354,221)(354,186){13}
//: {14}(355,268)(355,278)(375,278)(375,141){15}
output RegWrite;    //: /sn:0 /dp:1 {0}(680,221)(717,221)(717,220)(726,220){1}
output MemRead;    //: /sn:0 {0}(430,244)(414,244){1}
//: {2}(412,242)(412,221){3}
//: {4}(414,219)(424,219)(424,218)(659,218){5}
//: {6}(412,217)(412,119)(606,119){7}
//: {8}(610,119)(656,119){9}
//: {10}(608,121)(608,184)(658,184){11}
//: {12}(412,246)(412,274){13}
output MemToReg;    //: /sn:0 /dp:1 {0}(672,119)(714,119)(714,117)(724,117){1}
supply0 w5;    //: /sn:0 {0}(325,36)(408,36){1}
output Jump;    //: /sn:0 {0}(586,258)(564,258)(564,273){1}
wire w16;    //: /sn:0 {0}(254,336)(349,336){1}
//: {2}(353,336)(423,336){3}
//: {4}(427,336)(474,336){5}
//: {6}(478,336)(525,336){7}
//: {8}(529,336)(577,336)(577,294){9}
//: {10}(527,334)(527,294){11}
//: {12}(476,334)(476,295){13}
//: {14}(425,334)(425,295){15}
//: {16}(351,334)(351,296){17}
wire w6;    //: /sn:0 {0}(219,107)(241,107)(241,127)(263,127){1}
wire w22;    //: /sn:0 /dp:1 {0}(329,109)(329,167)(289,167){1}
wire w0;    //: /sn:0 /dp:1 {0}(373,101)(373,120){1}
wire w20;    //: /sn:0 {0}(376,80)(376,46)(408,46){1}
wire w12;    //: /sn:0 {0}(376,296)(376,375){1}
//: {2}(378,377)(398,377){3}
//: {4}(402,377)(449,377){5}
//: {6}(453,377)(500,377){7}
//: {8}(504,377)(552,377)(552,294){9}
//: {10}(502,375)(502,294){11}
//: {12}(451,375)(451,295){13}
//: {14}(400,375)(400,295){15}
//: {16}(374,377)(254,377){17}
wire w18;    //: /sn:0 {0}(219,164)(246,164){1}
//: {2}(250,164)(268,164){3}
//: {4}(248,166)(248,202)(349,202)(349,186){5}
wire w19;    //: /sn:0 {0}(219,187)(242,187)(242,169)(268,169){1}
wire w10;    //: /sn:0 {0}(567,294)(567,353)(519,353){1}
//: {2}(517,351)(517,294){3}
//: {4}(515,353)(468,353){5}
//: {6}(466,351)(466,295){7}
//: {8}(464,353)(417,353){9}
//: {10}(415,351)(415,295){11}
//: {12}(413,353)(363,353){13}
//: {14}(361,351)(361,296){15}
//: {16}(359,353)(254,353){17}
wire w23;    //: /sn:0 {0}(329,88)(329,66)(408,66){1}
wire w21;    //: /sn:0 /dp:1 {0}(324,109)(324,130)(284,130){1}
wire w8;    //: /sn:0 {0}(562,294)(562,361)(514,361){1}
//: {2}(512,359)(512,294){3}
//: {4}(510,361)(463,361){5}
//: {6}(461,359)(461,295){7}
//: {8}(459,361)(412,361){9}
//: {10}(410,359)(410,295){11}
//: {12}(408,361)(368,361){13}
//: {14}(366,359)(366,296){15}
//: {16}(364,361)(254,361){17}
wire w17;    //: /sn:0 {0}(352,165)(352,56)(408,56){1}
wire w14;    //: /sn:0 {0}(572,294)(572,345)(524,345){1}
//: {2}(522,343)(522,294){3}
//: {4}(520,345)(473,345){5}
//: {6}(471,343)(471,295){7}
//: {8}(469,345)(422,345){9}
//: {10}(420,343)(420,295){11}
//: {12}(418,345)(358,345){13}
//: {14}(356,343)(356,296){15}
//: {16}(354,345)(254,345){17}
wire w11;    //: /sn:0 {0}(371,296)(371,367){1}
//: {2}(373,369)(403,369){3}
//: {4}(407,369)(454,369){5}
//: {6}(458,369)(505,369){7}
//: {8}(509,369)(557,369)(557,294){9}
//: {10}(507,367)(507,294){11}
//: {12}(456,367)(456,295){13}
//: {14}(405,367)(405,295){15}
//: {16}(369,369)(254,369){17}
wire w15;    //: /sn:0 {0}(219,128)(225,128)(225,132)(248,132){1}
//: {2}(252,132)(263,132){3}
//: {4}(250,134)(250,150)(370,150)(370,141){5}
//: enddecls

  //: output g44 (Jump) @(583,258) /sn:0 /w:[ 0 ]
  nor g8 (.I0(w16), .I1(w14), .I2(w10), .I3(w8), .I4(w11), .I5(w12), .Z(RegDst));   //: @(363,285) /sn:0 /R:1 /w:[ 17 15 15 15 0 0 3 ]
  tran g4(.Z(w10), .I(Ins[28]));   //: @(248,353) /sn:0 /R:2 /w:[ 17 8 7 ] /ss:1
  or g75 (.I0(MemRead), .I1(RegDst), .Z(RegWrite));   //: @(670,221) /sn:0 /w:[ 5 11 0 ]
  //: output g47 (MemWrite) @(722,153) /sn:0 /w:[ 5 ]
  //: comment g16 /dolink:0 /link:"" @(398,279) /sn:0
  //: /line:"lw"
  //: /end
  tran g3(.Z(w14), .I(Ins[27]));   //: @(248,345) /sn:0 /R:2 /w:[ 17 6 5 ] /ss:1
  //: joint g26 (w12) @(451, 377) /w:[ 6 12 5 -1 ]
  and g17 (.I0(w12), .I1(!w11), .I2(w8), .I3(!w10), .I4(w14), .I5(w16), .Z(MemWrite));   //: @(463,284) /sn:0 /R:1 /w:[ 13 13 7 7 7 13 0 ]
  tran g2(.Z(w16), .I(Ins[26]));   //: @(248,336) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: joint g30 (w14) @(471, 345) /w:[ 5 6 8 -1 ]
  //: joint g23 (w16) @(425, 336) /w:[ 4 14 3 -1 ]
  //: joint g74 (MemWrite) @(558, 153) /w:[ 4 -1 3 6 ]
  //: comment g39 /dolink:0 /link:"" @(498,278) /sn:0
  //: /line:"beq"
  //: /end
  //: comment g24 /dolink:0 /link:"" @(449,280) /sn:0
  //: /line:"sw"
  //: /end
  //: comment g1 /dolink:0 /link:"" @(338,280) /sn:0
  //: /line:"Operacio"
  //: /end
  //: joint g77 (MemRead) @(412, 219) /w:[ 4 6 -1 3 ]
  //: joint g29 (w10) @(466, 353) /w:[ 5 6 8 -1 ]
  nand g60 (.I0(w18), .I1(RegDst), .Z(w17));   //: @(352,175) /sn:0 /R:1 /w:[ 5 13 0 ]
  //: joint g18 (w12) @(400, 377) /w:[ 4 14 3 -1 ]
  //: joint g70 (MemRead) @(412, 244) /w:[ 1 2 -1 12 ]
  and g25 (.I0(!w12), .I1(!w11), .I2(!w8), .I3(w10), .I4(!w14), .I5(!w16), .Z(Branch));   //: @(514,283) /sn:0 /R:1 /w:[ 11 11 3 3 3 11 5 ]
  //: joint g10 (w12) @(376, 377) /w:[ 2 1 16 -1 ]
  or g65 (.I0(w0), .I1(Branch), .Z(w20));   //: @(376,90) /sn:0 /R:1 /w:[ 0 0 0 ]
  //: joint g64 (w15) @(250, 132) /w:[ 2 -1 1 4 ]
  //: output g49 (RegWrite) @(723,220) /sn:0 /w:[ 1 ]
  or g72 (.I0(MemRead), .I1(MemWrite), .Z(ALUSrc));   //: @(669,187) /sn:0 /w:[ 11 7 0 ]
  concat g50 (.I0(w23), .I1(w17), .I2(w20), .I3(w5), .Z(ALUCtrl));   //: @(413,51) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  tran g6(.Z(w11), .I(Ins[30]));   //: @(248,369) /sn:0 /R:2 /w:[ 17 12 11 ] /ss:1
  //: joint g35 (w8) @(512, 361) /w:[ 1 2 4 -1 ]
  and g9 (.I0(w12), .I1(!w11), .I2(!w8), .I3(!w10), .I4(w14), .I5(w16), .Z(MemRead));   //: @(412,284) /sn:0 /R:1 /w:[ 15 15 11 11 11 15 13 ]
  tran g7(.Z(w12), .I(Ins[31]));   //: @(248,377) /sn:0 /R:2 /w:[ 17 14 13 ] /ss:1
  xor g56 (.I0(w18), .I1(w19), .Z(w22));   //: @(279,167) /sn:0 /w:[ 3 1 1 ]
  tran g58(.Z(w19), .I(Ins[3]));   //: @(213,187) /sn:0 /R:2 /w:[ 0 17 18 ] /ss:1
  //: joint g68 (RegDst) @(354, 244) /w:[ 6 8 -1 5 ]
  //: joint g73 (MemRead) @(608, 119) /w:[ 8 -1 7 10 ]
  //: joint g31 (w16) @(476, 336) /w:[ 6 12 5 -1 ]
  //: joint g22 (w14) @(420, 345) /w:[ 9 10 12 -1 ]
  and g59 (.I0(w21), .I1(w22), .I2(RegDst), .Z(w23));   //: @(329,98) /sn:0 /R:1 /w:[ 0 0 0 0 ]
  //: joint g71 (MemWrite) @(463, 269) /w:[ 2 8 -1 1 ]
  //: joint g67 (Branch) @(514, 263) /w:[ -1 2 1 4 ]
  //: output g45 (MemRead) @(427,244) /sn:0 /w:[ 0 ]
  //: output g41 (ALUCtrl) @(431,51) /sn:0 /w:[ 1 ]
  //: joint g36 (w10) @(517, 353) /w:[ 1 2 4 -1 ]
  //: joint g33 (w12) @(502, 377) /w:[ 8 10 7 -1 ]
  tran g54(.Z(w6), .I(Ins[0]));   //: @(213,107) /sn:0 /R:2 /w:[ 0 23 24 ] /ss:1
  //: joint g52 (Ins) @(215, 330) /w:[ 2 16 1 -1 ]
  //: output g42 (ALUSrc) @(723,185) /sn:0 /w:[ 1 ]
  //: comment g40 /dolink:0 /link:"" @(551,278) /sn:0
  //: /line:"j"
  //: /end
  buf g69 (.I(MemRead), .Z(MemToReg));   //: @(662,119) /sn:0 /w:[ 9 0 ]
  //: supply0 g66 (w5) @(319,36) /sn:0 /R:3 /w:[ 0 ]
  //: joint g12 (w8) @(366, 361) /w:[ 13 14 16 -1 ]
  //: output g46 (MemToReg) @(721,117) /sn:0 /w:[ 1 ]
  //: joint g34 (w11) @(507, 369) /w:[ 8 10 7 -1 ]
  //: joint g28 (w8) @(461, 361) /w:[ 5 6 8 -1 ]
  tran g57(.Z(w18), .I(Ins[2]));   //: @(213,164) /sn:0 /R:2 /w:[ 0 19 20 ] /ss:1
  //: joint g14 (w14) @(356, 345) /w:[ 13 14 16 -1 ]
  //: joint g11 (w11) @(371, 369) /w:[ 2 1 16 -1 ]
  tran g5(.Z(w8), .I(Ins[29]));   //: @(248,361) /sn:0 /R:2 /w:[ 17 10 9 ] /ss:1
  //: joint g21 (w10) @(415, 353) /w:[ 9 10 12 -1 ]
  //: joint g19 (w11) @(405, 369) /w:[ 4 14 3 -1 ]
  //: joint g61 (w18) @(248, 164) /w:[ 2 -1 1 4 ]
  and g32 (.I0(!w12), .I1(!w11), .I2(!w8), .I3(!w10), .I4(w14), .I5(!w16), .Z(Jump));   //: @(564,283) /sn:0 /R:1 /w:[ 9 9 0 0 0 9 1 ]
  //: joint g20 (w8) @(410, 361) /w:[ 9 10 12 -1 ]
  and g63 (.I0(w15), .I1(RegDst), .Z(w0));   //: @(373,130) /sn:0 /R:1 /w:[ 5 15 1 ]
  //: output g43 (Branch) @(532,254) /sn:0 /w:[ 3 ]
  //: joint g38 (w16) @(527, 336) /w:[ 8 10 7 -1 ]
  //: joint g15 (w16) @(351, 336) /w:[ 2 16 1 -1 ]
  //: input g0 (Ins) @(200,330) /sn:0 /w:[ 0 ]
  //: output g48 (RegDst) @(370,243) /sn:0 /w:[ 7 ]
  //: joint g27 (w11) @(456, 369) /w:[ 6 12 5 -1 ]
  //: joint g37 (w14) @(522, 345) /w:[ 1 2 4 -1 ]
  //: joint g62 (RegDst) @(355, 266) /w:[ 2 4 1 14 ]
  tran g55(.Z(w15), .I(Ins[1]));   //: @(213,128) /sn:0 /R:2 /w:[ 0 21 22 ] /ss:1
  //: joint g13 (w10) @(361, 353) /w:[ 13 14 16 -1 ]
  xor g53 (.I0(w6), .I1(w15), .Z(w21));   //: @(274,130) /sn:0 /w:[ 1 3 1 ]
  //: joint g76 (RegDst) @(354, 223) /w:[ 10 12 -1 9 ]

endmodule

module memoria(RD, WD, Addr, MemRead, MemWrite, clk);
//: interface  /sz:(297, 200) /bd:[ Ti0>MemWrite(147/297) Li0>WD[31:0](133/200) Li1>Addr[31:0](37/200) Bi0>clk(224/297) Bi1>MemRead(133/297) Ro0<RD[31:0](82/200) ]
supply0 w0;    //: /sn:0 {0}(715,297)(715,278){1}
input [31:0] Addr;    //: /sn:0 {0}(668,253)(704,253){1}
input [31:0] WD;    //: /sn:0 /dp:1 {0}(786,224)(786,201)(771,201){1}
input MemWrite;    //: /sn:0 {0}(623,163)(718,163){1}
//: {2}(722,163)(809,163)(809,232)(791,232){3}
//: {4}(720,165)(720,181){5}
input clk;    //: /sn:0 {0}(637,147)(725,147)(725,181){1}
output [31:0] RD;    //: /sn:0 {0}(833,251)(788,251){1}
//: {2}(786,249)(786,240){3}
//: {4}(784,251)(739,251){5}
input MemRead;    //: /sn:0 {0}(683,339)(729,339)(729,278){1}
wire w9;    //: /sn:0 {0}(722,202)(722,228){1}
//: enddecls

  //: output g4 (RD) @(830,251) /sn:0 /w:[ 0 ]
  bufif1 g8 (.Z(RD), .I(WD), .E(MemWrite));   //: @(786,230) /sn:0 /R:3 /w:[ 3 0 3 ]
  //: input g3 (WD) @(769,201) /sn:0 /w:[ 1 ]
  //: supply0 g2 (w0) @(715,303) /sn:0 /w:[ 0 ]
  //: input g1 (Addr) @(666,253) /sn:0 /w:[ 0 ]
  //: joint g10 (MemWrite) @(720, 163) /w:[ 2 -1 1 4 ]
  //: input g6 (MemRead) @(681,339) /sn:0 /w:[ 0 ]
  //: input g7 (MemWrite) @(621,163) /sn:0 /w:[ 0 ]
  nand g9 (.I0(clk), .I1(MemWrite), .Z(w9));   //: @(722,192) /sn:0 /R:3 /w:[ 1 5 0 ]
  //: joint g11 (RD) @(786, 251) /w:[ 1 2 4 -1 ]
  //: input g5 (clk) @(635,147) /sn:0 /w:[ 0 ]
  ram g0 (.A(Addr), .D(RD), .WE(w9), .OE(!MemRead), .CS(w0));   //: @(722,252) /sn:0 /w:[ 1 5 1 1 1 ]

endmodule

module ALU(AluOp, B, AluResult, Z, A);
//: interface  /sz:(40, 40) /bd:[ Ti0>op[3:0](20/40) Li0>a[31:0](10/40) Li1>b[31:0](30/40) Ro0<Q[31:0](30/40) Ro1<Z(10/40) ]
input [31:0] B;    //: /sn:0 {0}(-119,139)(-177,139)(-177,93){1}
//: {2}(-175,91)(-96,91)(-96,85)(-12,85){3}
//: {4}(-177,89)(-177,50)(-187,50){5}
input [31:0] A;    //: /sn:0 {0}(-202,-145)(-91,-145){1}
//: {2}(-87,-145)(92,-145){3}
//: {4}(96,-145)(119,-145)(119,-143)(136,-143){5}
//: {6}(94,-143)(94,-91)(143,-91){7}
//: {8}(-89,-143)(-89,-2)(157,-2){9}
output Z;    //: /sn:0 {0}(469,-32)(560,-32){1}
supply0 [30:0] w12;    //: /sn:0 {0}(217,51)(217,82)(237,82){1}
output [31:0] AluResult;    //: /sn:0 {0}(355,8)(394,8){1}
//: {2}(396,6)(396,-32)(448,-32){3}
//: {4}(396,10)(396,24)(543,24){5}
input [3:0] AluOp;    //: /sn:0 /dp:5 {0}(-174,204)(-21,204){1}
//: {2}(-20,204)(218,204){3}
//: {4}(219,204)(381,204){5}
wire [31:0] w7;    //: /sn:0 {0}(186,14)(199,14)(199,15)(205,15){1}
//: {2}(206,15)(270,15)(270,14)(326,14){3}
wire [1:0] w4;    //: /sn:0 {0}(219,199)(219,166)(342,166)(342,31){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(326,2)(296,2)(296,-93)(164,-93){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(157,30)(77,30)(77,75)(43,75){1}
//: {2}(41,73)(41,21){3}
//: {4}(43,19)(53,19)(53,-96)(143,-96){5}
//: {6}(41,17)(41,-138)(136,-138){7}
//: {8}(39,75)(17,75){9}
wire w1;    //: /sn:0 {0}(206,19)(206,92)(237,92){1}
wire w8;    //: /sn:0 {0}(-20,199)(-20,195)(4,195)(4,157){1}
//: {2}(6,155)(107,155)(107,-20)(171,-20)(171,-10){3}
//: {4}(4,153)(4,98){5}
wire [31:0] w14;    //: /sn:0 {0}(-103,139)(-57,139)(-57,65)(-12,65){1}
wire [31:0] w2;    //: /sn:0 {0}(157,-140)(316,-140)(316,-10)(326,-10){1}
wire w5;    //: /sn:0 /dp:1 {0}(172,79)(172,39)(171,39)(171,38){1}
wire [31:0] w9;    //: /sn:0 {0}(243,87)(319,87)(319,26)(326,26){1}
//: enddecls

  not g8 (.I(B), .Z(w14));   //: @(-113,139) /sn:0 /w:[ 0 0 ]
  or g4 (.I0(w0), .I1(A), .Z(w3));   //: @(154,-93) /sn:0 /w:[ 5 7 1 ]
  //: supply0 g16 (w12) @(217,45) /sn:0 /R:2 /w:[ 0 ]
  and g3 (.I0(A), .I1(w0), .Z(w2));   //: @(147,-140) /sn:0 /w:[ 5 7 0 ]
  tran g17(.Z(w1), .I(w7[31]));   //: @(206,13) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: input g2 (AluOp) @(-176,204) /sn:0 /w:[ 0 ]
  nor g23 (.I0(AluResult), .Z(Z));   //: @(459,-32) /sn:0 /w:[ 3 0 ]
  //: joint g24 (AluResult) @(396, 8) /w:[ -1 2 1 4 ]
  //: input g1 (B) @(-189,50) /sn:0 /w:[ 5 ]
  //: joint g18 (w8) @(4, 155) /w:[ 2 4 -1 1 ]
  //: joint g10 (A) @(-89, -145) /w:[ 2 -1 1 8 ]
  tran g6(.Z(w8), .I(AluOp[2]));   //: @(-20,202) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  add g9 (.A(w0), .B(A), .S(w7), .CI(w8), .CO(w5));   //: @(173,14) /sn:0 /R:1 /w:[ 0 9 0 3 1 ]
  //: joint g7 (B) @(-177, 91) /w:[ 2 4 -1 1 ]
  //: output g22 (AluResult) @(540,24) /sn:0 /w:[ 5 ]
  //: joint g12 (A) @(94, -145) /w:[ 4 -1 3 6 ]
  mux g14 (.I0(w2), .I1(w3), .I2(w7), .I3(w9), .S(w4), .Z(AluResult));   //: @(342,8) /sn:0 /R:1 /w:[ 1 0 3 1 1 0 ] /ss:0 /do:1
  //: joint g11 (w0) @(41, 75) /w:[ 1 2 8 -1 ]
  mux g5 (.I0(B), .I1(w14), .S(w8), .Z(w0));   //: @(4,75) /sn:0 /R:1 /w:[ 3 1 5 9 ] /ss:0 /do:0
  //: output g21 (Z) @(557,-32) /sn:0 /w:[ 1 ]
  led g19 (.I(w5));   //: @(172,86) /sn:0 /R:2 /w:[ 0 ] /type:0
  tran g20(.Z(w4), .I(AluOp[1:0]));   //: @(219,202) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:0
  concat g15 (.I0(w1), .I1(w12), .Z(w9));   //: @(242,87) /sn:0 /w:[ 1 1 0 ] /dr:0
  //: input g0 (A) @(-204,-145) /sn:0 /w:[ 0 ]
  //: joint g13 (w0) @(41, 19) /w:[ 4 6 -1 3 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Li0>Read1[4:0](32/182) Li1>Read2[4:0](72/182) Li2>Write[4:0](108/182) Li3>WriteData[31:0](148/182) Bi0>clk(108/147) Bi1>RegWrite(40/147) Ro0<Data1[31:0](47/182) Ro1<Data2[31:0](139/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,98){1}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,98){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,138){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [1:0] w10;    //: /sn:0 {0}(-140,148)(-140,432)(646,432){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-34){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-34)(-27,-23)(106,-23)(106,-10){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Fetch(Inst, Reset, Clk, PCIn, PCOut);
//: interface  /sz:(107, 96) /bd:[ Ti0>PCIn[31:0](76/107) Ti1>PCIn[31:0](76/107) Li0>Clk(65/96) Li1>Reset(22/96) Li2>Reset(22/96) Li3>Clk(65/96) To0<PCOut[31:0](28/107) To1<PCOut[31:0](28/107) Ro0<Inst[31:0](49/96) Ro1<Inst[31:0](49/96) ]
supply0 w13;    //: /sn:0 {0}(348,222)(348,195){1}
output [31:0] PCOut;    //: /sn:0 /dp:1 {0}(429,76)(482,76){1}
input Clk;    //: /sn:0 {0}(188,208)(238,208)(238,185){1}
output [31:0] Inst;    //: /sn:0 {0}(427,168)(365,168){1}
input [31:0] PCIn;    //: /sn:0 {0}(148,147)(227,147){1}
input Reset;    //: /sn:0 {0}(182,91)(233,91)(233,109){1}
supply0 w14;    //: /sn:0 {0}(243,66)(243,109){1}
supply0 w15;    //: /sn:0 {0}(439,39)(414,39)(414,52){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(352,46)(352,60)(400,60){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(248,147)(301,147){1}
//: {2}(305,147)(326,147)(326,170)(330,170){3}
//: {4}(303,145)(303,92)(400,92){5}
wire w12;    //: /sn:0 {0}(414,100)(414,110){1}
//: enddecls

  //: output g8 (Inst) @(424,168) /sn:0 /w:[ 0 ]
  //: supply0 g4 (w14) @(243,60) /sn:0 /R:2 /w:[ 0 ]
  //: supply0 g3 (w13) @(348,228) /sn:0 /w:[ 0 ]
  add g2 (.A(w3), .B(w0), .S(PCOut), .CI(w15), .CO(w12));   //: @(416,76) /sn:0 /R:1 /w:[ 5 1 0 1 0 ]
  register g1 (.Q(w3), .D(PCIn), .EN(w14), .CLR(!Reset), .CK(!Clk));   //: @(238,147) /sn:0 /R:1 /w:[ 0 1 1 1 1 ]
  //: input g10 (Reset) @(180,91) /sn:0 /w:[ 0 ]
  //: joint g6 (w3) @(303, 147) /w:[ 2 4 1 -1 ]
  //: input g9 (Clk) @(186,208) /sn:0 /w:[ 0 ]
  //: dip g7 (w0) @(352,36) /sn:0 /w:[ 0 ] /st:1
  //: input g12 (PCIn) @(146,147) /sn:0 /w:[ 0 ]
  //: output g11 (PCOut) @(479,76) /sn:0 /w:[ 1 ]
  //: supply0 g5 (w15) @(445,39) /sn:0 /R:1 /w:[ 0 ]
  rom g0 (.A(w3), .D(Inst), .OE(w13));   //: @(348,169) /sn:0 /w:[ 3 1 1 ] /mem:"/media/sf_Carpeta_Compartida_Linux/EC-2/mult.mem"

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clk, clr, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Li0>clk(59/69) Li1>RegWr(47/69) Li2>SB[2:0](22/69) Li3>SA[2:0](11/69) Li4>SD[2:0](35/69) Ri0>clr(35/69) Bo0<BOUT[31:0](65/98) Bo1<AOUT[31:0](37/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module Read(SignExOut, SignExIn, RegDst, R1, R2, WR, RD2, RD1, WriteData, clk, clr, RegWrite);
//: interface  /sz:(162, 244) /bd:[ Ti0>RegWrite(85/162) Ti1>RegWrite(85/162) Li0>SignExIn[15:0](200/244) Li1>WriteData[31:0](153/244) Li2>RegDst(122/244) Li3>WR[4:0](97/244) Li4>R2[4:0](65/244) Li5>R1[4:0](34/244) Li6>SignExIn[15:0](200/244) Li7>WriteData[31:0](153/244) Li8>RegDst(122/244) Li9>WR[4:0](97/244) Li10>R2[4:0](65/244) Li11>R1[4:0](34/244) Bi0>clr(111/162) Bi1>clk(55/162) Bi2>clr(111/162) Bi3>clk(55/162) Ro0<SignExOut[31:0](205/244) Ro1<RD2[31:0](126/244) Ro2<RD1[31:0](49/244) Ro3<SignExOut[31:0](205/244) Ro4<RD2[31:0](126/244) Ro5<RD1[31:0](49/244) ]
input [4:0] WR;    //: /sn:0 /dp:1 {0}(480,219)(411,219){1}
input [4:0] R2;    //: /sn:0 {0}(412,173)(439,173){1}
//: {2}(443,173)(532,173){3}
//: {4}(441,175)(441,199)(480,199){5}
input [31:0] WriteData;    //: /sn:0 {0}(407,249)(532,249){1}
output [31:0] SignExOut;    //: /sn:0 {0}(718,440)(637,440){1}
output [31:0] RD2;    //: /sn:0 {0}(720,240)(681,240){1}
input [4:0] R1;    //: /sn:0 {0}(411,133)(532,133){1}
input RegDst;    //: /sn:0 {0}(448,332)(471,332)(471,176)(496,176)(496,186){1}
input clr;    //: /sn:0 {0}(585,65)(599,65)(599,100){1}
input RegWrite;    //: /sn:0 {0}(565,324)(573,324)(573,284){1}
input clk;    //: /sn:0 {0}(624,322)(641,322)(641,284){1}
output [31:0] RD1;    //: /sn:0 {0}(724,148)(681,148){1}
input [15:0] SignExIn;    //: /sn:0 {0}(499,441)(571,441){1}
wire [4:0] w12;    //: /sn:0 /dp:1 {0}(509,209)(532,209){1}
//: enddecls

  //: output g4 (SignExOut) @(715,440) /sn:0 /w:[ 0 ]
  //: joint g8 (R2) @(441, 173) /w:[ 2 -1 1 4 ]
  //: input g3 (SignExIn) @(497,441) /sn:0 /w:[ 0 ]
  mux g2 (.I0(R2), .I1(WR), .S(RegDst), .Z(w12));   //: @(496,209) /sn:0 /R:1 /w:[ 5 0 1 0 ] /ss:1 /do:1
  Sign_extend g1 (.in(SignExIn), .out(SignExOut));   //: @(572, 404) /sz:(64, 66) /sn:0 /p:[ Li0>1 Ro0<1 ]
  //: input g10 (RegDst) @(446,332) /sn:0 /w:[ 0 ]
  //: input g6 (R1) @(409,133) /sn:0 /w:[ 0 ]
  //: input g7 (R2) @(410,173) /sn:0 /w:[ 0 ]
  //: input g9 (WR) @(409,219) /sn:0 /w:[ 1 ]
  //: output g12 (RD2) @(717,240) /sn:0 /w:[ 0 ]
  //: output g11 (RD1) @(721,148) /sn:0 /w:[ 0 ]
  //: input g5 (WriteData) @(405,249) /sn:0 /w:[ 0 ]
  //: input g14 (clk) @(622,322) /sn:0 /w:[ 0 ]
  //: input g15 (clr) @(583,65) /sn:0 /w:[ 0 ]
  BRegs32x32 g0 (.clr(clr), .Read1(R1), .Read2(R2), .Write(w12), .WriteData(WriteData), .clk(clk), .RegWrite(RegWrite), .Data1(RD1), .Data2(RD2));   //: @(533, 101) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>1 Li1>3 Li2>1 Li3>1 Bi0>1 Bi1>1 Ro0<1 Ro1<1 ]
  //: input g13 (RegWrite) @(563,324) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [4:0] w16;    //: /sn:0 {0}(548,200)(485,200){1}
wire [31:0] w13;    //: /sn:0 {0}(956,271)(977,271){1}
//: {2}(981,271)(991,271)(991,270)(1001,270){3}
//: {4}(979,269)(979,246)(989,246)(989,198)(1143,198)(1143,180){5}
//: {6}(979,273)(979,400)(1211,400)(1211,319)(1256,319){7}
wire w34;    //: /sn:0 /dp:1 {0}(808,13)(808,-87)(314,-87){1}
wire [25:0] w4;    //: /sn:0 {0}(733,33)(485,33){1}
wire [31:0] w25;    //: /sn:0 {0}(712,340)(771,340)(771,283){1}
//: {2}(773,281)(801,281){3}
//: {4}(771,279)(771,95){5}
wire [31:0] w0;    //: /sn:0 {0}(393,351)(393,-21)(879,-21)(879,28){1}
//: {2}(881,30)(1054,30)(1054,22){3}
//: {4}(879,32)(879,50)(856,50){5}
wire w36;    //: /sn:0 /dp:1 {0}(1272,286)(1272,-46)(314,-46){1}
wire [31:0] w22;    //: /sn:0 /dp:1 {0}(830,271)(884,271){1}
wire [15:0] w20;    //: /sn:0 {0}(548,335)(485,335){1}
wire w42;    //: /sn:0 {0}(821,134)(821,172)(974,172)(974,239)(956,239){1}
wire w19;    //: /sn:0 {0}(314,-8)(1094,-8)(1094,247){1}
wire [3:0] w18;    //: /sn:0 /dp:1 {0}(314,-26)(920,-26)(920,222){1}
wire [31:0] w23;    //: /sn:0 /dp:1 {0}(1256,299)(1199,299)(1199,298)(1189,298){1}
wire w10;    //: /sn:0 /dp:1 {0}(816,134)(816,147)(848,147)(848,-111)(314,-111){1}
wire w21;    //: /sn:0 {0}(314,10)(726,10)(726,206)(802,206)(802,238)(817,238)(817,248){1}
wire [31:0] w24;    //: /sn:0 {0}(1001,329)(743,329)(743,263){1}
//: {2}(745,261)(778,261){3}
//: {4}(782,261)(801,261){5}
//: {6}(780,263)(780,386){7}
//: {8}(741,261)(712,261){9}
wire [31:0] w1;    //: /sn:0 {0}(180,-59)(152,-59)(152,122)(480,122){1}
//: {2}(482,120)(482,33){3}
//: {4}(482,32)(482,25){5}
//: {6}(482,124)(482,168){7}
//: {8}(482,169)(482,199){9}
//: {10}(482,200)(482,231){11}
//: {12}(482,232)(482,295){13}
//: {14}(480,297)(207,297)(207,257){15}
//: {16}(482,299)(482,334){17}
//: {18}(482,335)(482,401)(425,401){19}
wire [31:0] w31;    //: /sn:0 /dp:1 {0}(1285,309)(1293,309)(1293,366){1}
//: {2}(1295,368)(1421,368)(1421,342){3}
//: {4}(1293,370)(1293,433)(534,433)(534,288)(548,288){5}
wire w32;    //: /sn:0 /dp:1 {0}(548,257)(506,257)(506,-133)(314,-133){1}
wire [4:0] w17;    //: /sn:0 {0}(548,232)(485,232){1}
wire w27;    //: /sn:0 {0}(134,569)(272,569){1}
//: {2}(276,569)(602,569){3}
//: {4}(606,569)(1142,569)(1142,371){5}
//: {6}(604,567)(604,380){7}
//: {8}(274,567)(274,417)(316,417){9}
wire w28;    //: /sn:0 {0}(314,28)(613,28)(613,108)(634,108)(634,134){1}
wire w35;    //: /sn:0 /dp:1 {0}(1085,371)(1085,459)(1530,459)(1530,-68)(314,-68){1}
wire w2;    //: /sn:0 {0}(223,375)(284,375){1}
//: {2}(288,375)(302,375)(302,374)(316,374){3}
//: {4}(286,377)(286,483)(660,483)(660,380){5}
wire [31:0] w11;    //: /sn:0 {0}(884,239)(843,239)(843,186){1}
//: {2}(845,184)(1001,184)(1001,127){3}
//: {4}(841,184)(712,184){5}
wire [4:0] w15;    //: /sn:0 {0}(548,169)(485,169){1}
wire w43;    //: /sn:0 {0}(819,113)(819,95){1}
wire [31:0] w26;    //: /sn:0 {0}(345,351)(345,65)(733,65){1}
//: enddecls

  clock g4 (.Z(w27));   //: @(121,569) /sn:0 /w:[ 0 ] /omega:2000 /phi:0 /duty:50
  tran g8(.Z(w15), .I(w1[25:21]));   //: @(480,169) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  UC g16 (.Ins(w1), .RegWrite(w28), .ALUSrc(w21), .MemWrite(w19), .ALUCtrl(w18), .MemToReg(w36), .MemRead(w35), .Jump(w34), .Branch(w10), .RegDst(w32));   //: @(181, -155) /sz:(132, 211) /sn:0 /p:[ Li0>0 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<1 Ro5<1 Ro6<1 Ro7<1 Ro8<1 ]
  Read g3 (.RegWrite(w28), .SignExIn(w20), .WriteData(w31), .RegDst(w32), .WR(w17), .R2(w16), .R1(w15), .clr(w2), .clk(w27), .SignExOut(w25), .RD2(w24), .RD1(w11));   //: @(549, 135) /sz:(162, 244) /sn:0 /p:[ Ti0>1 Li0>0 Li1>5 Li2>0 Li3>0 Li4>0 Li5>0 Bi0>5 Bi1>7 Ro0<0 Ro1<9 Ro2<5 ]
  //: joint g17 (w1) @(482, 122) /w:[ -1 2 1 6 ]
  ALU g2 (.AluOp(w18), .A(w11), .B(w22), .AluResult(w13), .Z(w42));   //: @(885, 223) /sz:(70, 65) /sn:0 /p:[ Ti0>1 Li0>0 Li1>1 Ro0<0 Ro1<1 ]
  //: joint g23 (w13) @(979, 271) /w:[ 2 4 1 6 ]
  led g30 (.I(w0));   //: @(1054,15) /sn:0 /w:[ 3 ] /type:2
  jump g1 (.jump(w34), .PCNext(w26), .inm26(w4), .PCSrc(w43), .SignXtended(w25), .dir(w0));   //: @(734, 14) /sz:(121, 80) /sn:0 /p:[ Ti0>0 Li0>1 Li1>0 Bi0>1 Bi1>5 Ro0<5 ]
  //: joint g39 (w24) @(780, 261) /w:[ 4 -1 3 6 ]
  //: joint g29 (w31) @(1293, 368) /w:[ 2 1 -1 4 ]
  tran g10(.Z(w17), .I(w1[15:11]));   //: @(480,232) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  //: switch g6 (w2) @(206,375) /sn:0 /w:[ 0 ] /st:0
  //: joint g7 (w2) @(286, 375) /w:[ 2 -1 1 4 ]
  tran g9(.Z(w16), .I(w1[20:16]));   //: @(480,200) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  //: joint g31 (w0) @(879, 30) /w:[ 2 1 -1 4 ]
  //: joint g22 (w27) @(604, 569) /w:[ 4 6 3 -1 ]
  led g36 (.I(w11));   //: @(1001,120) /sn:0 /w:[ 3 ] /type:2
  //: joint g33 (w1) @(482, 297) /w:[ -1 13 14 16 ]
  led g40 (.I(w13));   //: @(1143,173) /sn:0 /w:[ 5 ] /type:2
  tran g12(.Z(w4), .I(w1[25:0]));   //: @(480,33) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  led g28 (.I(w31));   //: @(1421,335) /sn:0 /w:[ 3 ] /type:2
  //: joint g5 (w27) @(274, 569) /w:[ 2 8 1 -1 ]
  tran g11(.Z(w20), .I(w1[15:0]));   //: @(480,335) /sn:0 /R:2 /w:[ 1 18 17 ] /ss:1
  //: joint g14 (w25) @(771, 281) /w:[ 2 4 -1 1 ]
  memoria g19 (.MemWrite(w19), .WD(w24), .Addr(w13), .clk(w27), .MemRead(w35), .RD(w23));   //: @(1002, 248) /sz:(186, 122) /sn:0 /p:[ Ti0>1 Li0>0 Li1>3 Bi0>5 Bi1>0 Ro0<1 ]
  mux g21 (.I0(w13), .I1(w23), .S(w36), .Z(w31));   //: @(1272,309) /sn:0 /R:1 /w:[ 7 0 0 0 ] /ss:1 /do:1
  led g32 (.I(w1));   //: @(207,250) /sn:0 /w:[ 15 ] /type:2
  //: joint g20 (w24) @(743, 261) /w:[ 2 -1 8 1 ]
  led g38 (.I(w24));   //: @(780,393) /sn:0 /R:2 /w:[ 7 ] /type:2
  and g15 (.I0(w10), .I1(w42), .Z(w43));   //: @(819,123) /sn:0 /R:1 /w:[ 0 0 0 ]
  Fetch g0 (.PCIn(w0), .Reset(w2), .Clk(w27), .PCOut(w26), .Inst(w1));   //: @(317, 352) /sz:(107, 96) /sn:0 /p:[ Ti0>0 Li0>3 Li1>9 To0<0 Ro0<19 ]
  //: joint g37 (w11) @(843, 184) /w:[ 2 -1 4 1 ]
  mux g13 (.I0(w24), .I1(w25), .S(w21), .Z(w22));   //: @(817,271) /sn:0 /R:1 /w:[ 5 3 1 0 ] /ss:1 /do:1

endmodule

module Sign_extend(out, in);
//: interface  /sz:(64, 66) /bd:[ Li0>in[15:0](37/66) Ro0<out[31:0](36/66) ]
input [15:0] in;    //: /sn:0 {0}(441,165)(464,165)(464,166){1}
//: {2}(464,167)(464,350){3}
//: {4}(464,351)(464,359){5}
output [31:0] out;    //: /sn:0 {0}(606,266)(571,266){1}
wire [14:0] w0;    //: /sn:0 {0}(467,351)(565,351){1}
wire w18;    //: /sn:0 {0}(565,181)(473,181){1}
//: {2}(471,179)(471,167)(467,167){3}
//: {4}(471,183)(471,199){5}
//: {6}(473,201)(521,201){7}
//: {8}(525,201)(565,201){9}
//: {10}(523,199)(523,191)(565,191){11}
//: {12}(471,203)(471,219){13}
//: {14}(473,221)(521,221){15}
//: {16}(525,221)(565,221){17}
//: {18}(523,219)(523,211)(565,211){19}
//: {20}(471,223)(471,239){21}
//: {22}(473,241)(521,241){23}
//: {24}(525,241)(565,241){25}
//: {26}(523,239)(523,231)(565,231){27}
//: {28}(471,243)(471,259){29}
//: {30}(473,261)(521,261){31}
//: {32}(525,261)(565,261){33}
//: {34}(523,259)(523,251)(565,251){35}
//: {36}(471,263)(471,279){37}
//: {38}(473,281)(520,281){39}
//: {40}(524,281)(565,281){41}
//: {42}(522,279)(522,271)(565,271){43}
//: {44}(471,283)(471,299){45}
//: {46}(473,301)(520,301){47}
//: {48}(524,301)(565,301){49}
//: {50}(522,299)(522,291)(565,291){51}
//: {52}(471,303)(471,319){53}
//: {54}(473,321)(519,321){55}
//: {56}(523,321)(565,321){57}
//: {58}(521,319)(521,311)(565,311){59}
//: {60}(471,323)(471,339){61}
//: {62}(473,341)(519,341){63}
//: {64}(523,341)(565,341){65}
//: {66}(521,339)(521,331)(565,331){67}
//: {68}(471,343)(471,348){69}
//: enddecls

  tran g4(.Z(w18), .I(in[15]));   //: @(462,167) /sn:0 /R:2 /w:[ 3 2 1 ] /ss:1
  //: joint g8 (w18) @(521, 321) /w:[ 56 58 55 -1 ]
  tran g3(.Z(w0), .I(in[14:0]));   //: @(462,351) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: joint g16 (w18) @(523, 241) /w:[ 24 26 23 -1 ]
  //: joint g17 (w18) @(471, 221) /w:[ 14 13 -1 20 ]
  concat g2 (.I0(w0), .I1(w18), .I2(w18), .I3(w18), .I4(w18), .I5(w18), .I6(w18), .I7(w18), .I8(w18), .I9(w18), .I10(w18), .I11(w18), .I12(w18), .I13(w18), .I14(w18), .I15(w18), .I16(w18), .I17(w18), .Z(out));   //: @(570,266) /sn:0 /w:[ 1 65 67 57 59 49 51 41 43 33 35 25 27 17 19 9 11 0 1 ] /dr:0
  //: output g1 (out) @(603,266) /sn:0 /w:[ 0 ]
  //: joint g18 (w18) @(523, 221) /w:[ 16 18 15 -1 ]
  //: joint g10 (w18) @(522, 301) /w:[ 48 50 47 -1 ]
  //: joint g6 (w18) @(521, 341) /w:[ 64 66 63 -1 ]
  //: joint g7 (w18) @(471, 321) /w:[ 54 53 -1 60 ]
  //: joint g9 (w18) @(471, 301) /w:[ 46 45 -1 52 ]
  //: joint g12 (w18) @(522, 281) /w:[ 40 42 39 -1 ]
  //: joint g11 (w18) @(471, 281) /w:[ 38 37 -1 44 ]
  //: joint g5 (w18) @(471, 341) /w:[ 62 61 -1 68 ]
  //: joint g14 (w18) @(523, 261) /w:[ 32 34 31 -1 ]
  //: joint g19 (w18) @(471, 201) /w:[ 6 5 -1 12 ]
  //: joint g21 (w18) @(471, 181) /w:[ 1 2 -1 4 ]
  //: joint g20 (w18) @(523, 201) /w:[ 8 10 7 -1 ]
  //: joint g15 (w18) @(471, 241) /w:[ 22 21 -1 28 ]
  //: input g0 (in) @(439,165) /sn:0 /w:[ 0 ]
  //: joint g13 (w18) @(471, 261) /w:[ 30 29 -1 36 ]

endmodule
